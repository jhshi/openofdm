///////////////////////////////////////////////////////////
//  Copyright (c) 1995/2006 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /    Vendor      : Xilinx 
// \  \    \/     Version : 10.1
//  \  \          Description : 
//  /  /                      
// /__/   /\      Filename    : PPC440.v
// \  \  /  \     Timestamp   : Thu Apr 19 10:07:12 2007

//  \__\/\__ \                    
//                                 
//  Generated by : SmartModelVerilogFileWriter (sm_verilog)
//  Revision:
///////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module PPC440 (
	APUFCMDECFPUOP,
	APUFCMDECLDSTXFERSIZE,
	APUFCMDECLOAD,
	APUFCMDECNONAUTON,
	APUFCMDECSTORE,
	APUFCMDECUDI,
	APUFCMDECUDIVALID,
	APUFCMENDIAN,
	APUFCMFLUSH,
	APUFCMINSTRUCTION,
	APUFCMINSTRVALID,
	APUFCMLOADBYTEADDR,
	APUFCMLOADDATA,
	APUFCMLOADDVALID,
	APUFCMMSRFE0,
	APUFCMMSRFE1,
	APUFCMNEXTINSTRREADY,
	APUFCMOPERANDVALID,
	APUFCMRADATA,
	APUFCMRBDATA,
	APUFCMWRITEBACKOK,
	C440CPMCORESLEEPREQ,
	C440CPMDECIRPTREQ,
	C440CPMFITIRPTREQ,
	C440CPMMSRCE,
	C440CPMMSREE,
	C440CPMTIMERRESETREQ,
	C440CPMWDIRPTREQ,
	C440DBGSYSTEMCONTROL,
	C440JTGTDO,
	C440JTGTDOEN,
	C440MACHINECHECK,
	C440RSTCHIPRESETREQ,
	C440RSTCORERESETREQ,
	C440RSTSYSTEMRESETREQ,
	C440TRCBRANCHSTATUS,
	C440TRCCYCLE,
	C440TRCEXECUTIONSTATUS,
	C440TRCTRACESTATUS,
	C440TRCTRIGGEREVENTOUT,
	C440TRCTRIGGEREVENTTYPE,
	DMA0LLRSTENGINEACK,
	DMA0LLRXDSTRDYN,
	DMA0LLTXD,
	DMA0LLTXEOFN,
	DMA0LLTXEOPN,
	DMA0LLTXREM,
	DMA0LLTXSOFN,
	DMA0LLTXSOPN,
	DMA0LLTXSRCRDYN,
	DMA0RXIRQ,
	DMA0TXIRQ,
	DMA1LLRSTENGINEACK,
	DMA1LLRXDSTRDYN,
	DMA1LLTXD,
	DMA1LLTXEOFN,
	DMA1LLTXEOPN,
	DMA1LLTXREM,
	DMA1LLTXSOFN,
	DMA1LLTXSOPN,
	DMA1LLTXSRCRDYN,
	DMA1RXIRQ,
	DMA1TXIRQ,
	DMA2LLRSTENGINEACK,
	DMA2LLRXDSTRDYN,
	DMA2LLTXD,
	DMA2LLTXEOFN,
	DMA2LLTXEOPN,
	DMA2LLTXREM,
	DMA2LLTXSOFN,
	DMA2LLTXSOPN,
	DMA2LLTXSRCRDYN,
	DMA2RXIRQ,
	DMA2TXIRQ,
	DMA3LLRSTENGINEACK,
	DMA3LLRXDSTRDYN,
	DMA3LLTXD,
	DMA3LLTXEOFN,
	DMA3LLTXEOPN,
	DMA3LLTXREM,
	DMA3LLTXSOFN,
	DMA3LLTXSOPN,
	DMA3LLTXSRCRDYN,
	DMA3RXIRQ,
	DMA3TXIRQ,
	MIMCADDRESS,
	MIMCADDRESSVALID,
	MIMCBANKCONFLICT,
	MIMCBYTEENABLE,
	MIMCREADNOTWRITE,
	MIMCROWCONFLICT,
	MIMCWRITEDATA,
	MIMCWRITEDATAVALID,
	PPCCPMINTERCONNECTBUSY,
	PPCDMDCRABUS,
	PPCDMDCRDBUSOUT,
	PPCDMDCRREAD,
	PPCDMDCRUABUS,
	PPCDMDCRWRITE,
	PPCDSDCRACK,
	PPCDSDCRDBUSIN,
	PPCDSDCRTIMEOUTWAIT,
	PPCEICINTERCONNECTIRQ,
	PPCMPLBABORT,
	PPCMPLBABUS,
	PPCMPLBBE,
	PPCMPLBBUSLOCK,
	PPCMPLBLOCKERR,
	PPCMPLBPRIORITY,
	PPCMPLBRDBURST,
	PPCMPLBREQUEST,
	PPCMPLBRNW,
	PPCMPLBSIZE,
	PPCMPLBTATTRIBUTE,
	PPCMPLBTYPE,
	PPCMPLBUABUS,
	PPCMPLBWRBURST,
	PPCMPLBWRDBUS,
	PPCS0PLBADDRACK,
	PPCS0PLBMBUSY,
	PPCS0PLBMIRQ,
	PPCS0PLBMRDERR,
	PPCS0PLBMWRERR,
	PPCS0PLBRDBTERM,
	PPCS0PLBRDCOMP,
	PPCS0PLBRDDACK,
	PPCS0PLBRDDBUS,
	PPCS0PLBRDWDADDR,
	PPCS0PLBREARBITRATE,
	PPCS0PLBSSIZE,
	PPCS0PLBWAIT,
	PPCS0PLBWRBTERM,
	PPCS0PLBWRCOMP,
	PPCS0PLBWRDACK,
	PPCS1PLBADDRACK,
	PPCS1PLBMBUSY,
	PPCS1PLBMIRQ,
	PPCS1PLBMRDERR,
	PPCS1PLBMWRERR,
	PPCS1PLBRDBTERM,
	PPCS1PLBRDCOMP,
	PPCS1PLBRDDACK,
	PPCS1PLBRDDBUS,
	PPCS1PLBRDWDADDR,
	PPCS1PLBREARBITRATE,
	PPCS1PLBSSIZE,
	PPCS1PLBWAIT,
	PPCS1PLBWRBTERM,
	PPCS1PLBWRCOMP,
	PPCS1PLBWRDACK,

	CPMC440CLK,
	CPMC440CLKEN,
	CPMC440CORECLOCKINACTIVE,
	CPMC440TIMERCLOCK,
	CPMDCRCLK,
	CPMDMA0LLCLK,
	CPMDMA1LLCLK,
	CPMDMA2LLCLK,
	CPMDMA3LLCLK,
	CPMFCMCLK,
	CPMINTERCONNECTCLK,
	CPMINTERCONNECTCLKEN,
	CPMINTERCONNECTCLKNTO1,
	CPMMCCLK,
	CPMPPCMPLBCLK,
	CPMPPCS0PLBCLK,
	CPMPPCS1PLBCLK,
	DBGC440DEBUGHALT,
	DBGC440SYSTEMSTATUS,
	DBGC440UNCONDDEBUGEVENT,
	DCRPPCDMACK,
	DCRPPCDMDBUSIN,
	DCRPPCDMTIMEOUTWAIT,
	DCRPPCDSABUS,
	DCRPPCDSDBUSOUT,
	DCRPPCDSREAD,
	DCRPPCDSWRITE,
	EICC440CRITIRQ,
	EICC440EXTIRQ,
	FCMAPUCONFIRMINSTR,
	FCMAPUCR,
	FCMAPUDONE,
	FCMAPUEXCEPTION,
	FCMAPUFPSCRFEX,
	FCMAPURESULT,
	FCMAPURESULTVALID,
	FCMAPUSLEEPNOTREADY,
	FCMAPUSTOREDATA,
	JTGC440TCK,
	JTGC440TDI,
	JTGC440TMS,
	JTGC440TRSTNEG,
	LLDMA0RSTENGINEREQ,
	LLDMA0RXD,
	LLDMA0RXEOFN,
	LLDMA0RXEOPN,
	LLDMA0RXREM,
	LLDMA0RXSOFN,
	LLDMA0RXSOPN,
	LLDMA0RXSRCRDYN,
	LLDMA0TXDSTRDYN,
	LLDMA1RSTENGINEREQ,
	LLDMA1RXD,
	LLDMA1RXEOFN,
	LLDMA1RXEOPN,
	LLDMA1RXREM,
	LLDMA1RXSOFN,
	LLDMA1RXSOPN,
	LLDMA1RXSRCRDYN,
	LLDMA1TXDSTRDYN,
	LLDMA2RSTENGINEREQ,
	LLDMA2RXD,
	LLDMA2RXEOFN,
	LLDMA2RXEOPN,
	LLDMA2RXREM,
	LLDMA2RXSOFN,
	LLDMA2RXSOPN,
	LLDMA2RXSRCRDYN,
	LLDMA2TXDSTRDYN,
	LLDMA3RSTENGINEREQ,
	LLDMA3RXD,
	LLDMA3RXEOFN,
	LLDMA3RXEOPN,
	LLDMA3RXREM,
	LLDMA3RXSOFN,
	LLDMA3RXSOPN,
	LLDMA3RXSRCRDYN,
	LLDMA3TXDSTRDYN,
	MCMIADDRREADYTOACCEPT,
	MCMIREADDATA,
	MCMIREADDATAERR,
	MCMIREADDATAVALID,
	PLBPPCMADDRACK,
	PLBPPCMMBUSY,
	PLBPPCMMIRQ,
	PLBPPCMMRDERR,
	PLBPPCMMWRERR,
	PLBPPCMRDBTERM,
	PLBPPCMRDDACK,
	PLBPPCMRDDBUS,
	PLBPPCMRDPENDPRI,
	PLBPPCMRDPENDREQ,
	PLBPPCMRDWDADDR,
	PLBPPCMREARBITRATE,
	PLBPPCMREQPRI,
	PLBPPCMSSIZE,
	PLBPPCMTIMEOUT,
	PLBPPCMWRBTERM,
	PLBPPCMWRDACK,
	PLBPPCMWRPENDPRI,
	PLBPPCMWRPENDREQ,
	PLBPPCS0ABORT,
	PLBPPCS0ABUS,
	PLBPPCS0BE,
	PLBPPCS0BUSLOCK,
	PLBPPCS0LOCKERR,
	PLBPPCS0MASTERID,
	PLBPPCS0MSIZE,
	PLBPPCS0PAVALID,
	PLBPPCS0RDBURST,
	PLBPPCS0RDPENDPRI,
	PLBPPCS0RDPENDREQ,
	PLBPPCS0RDPRIM,
	PLBPPCS0REQPRI,
	PLBPPCS0RNW,
	PLBPPCS0SAVALID,
	PLBPPCS0SIZE,
	PLBPPCS0TATTRIBUTE,
	PLBPPCS0TYPE,
	PLBPPCS0UABUS,
	PLBPPCS0WRBURST,
	PLBPPCS0WRDBUS,
	PLBPPCS0WRPENDPRI,
	PLBPPCS0WRPENDREQ,
	PLBPPCS0WRPRIM,
	PLBPPCS1ABORT,
	PLBPPCS1ABUS,
	PLBPPCS1BE,
	PLBPPCS1BUSLOCK,
	PLBPPCS1LOCKERR,
	PLBPPCS1MASTERID,
	PLBPPCS1MSIZE,
	PLBPPCS1PAVALID,
	PLBPPCS1RDBURST,
	PLBPPCS1RDPENDPRI,
	PLBPPCS1RDPENDREQ,
	PLBPPCS1RDPRIM,
	PLBPPCS1REQPRI,
	PLBPPCS1RNW,
	PLBPPCS1SAVALID,
	PLBPPCS1SIZE,
	PLBPPCS1TATTRIBUTE,
	PLBPPCS1TYPE,
	PLBPPCS1UABUS,
	PLBPPCS1WRBURST,
	PLBPPCS1WRDBUS,
	PLBPPCS1WRPENDPRI,
	PLBPPCS1WRPENDREQ,
	PLBPPCS1WRPRIM,
	RSTC440RESETCHIP,
	RSTC440RESETCORE,
	RSTC440RESETSYSTEM,
	TIEC440DCURDLDCACHEPLBPRIO,
	TIEC440DCURDNONCACHEPLBPRIO,
	TIEC440DCURDTOUCHPLBPRIO,
	TIEC440DCURDURGENTPLBPRIO,
	TIEC440DCUWRFLUSHPLBPRIO,
	TIEC440DCUWRSTOREPLBPRIO,
	TIEC440DCUWRURGENTPLBPRIO,
	TIEC440ENDIANRESET,
	TIEC440ERPNRESET,
	TIEC440ICURDFETCHPLBPRIO,
	TIEC440ICURDSPECPLBPRIO,
	TIEC440ICURDTOUCHPLBPRIO,
	TIEC440PIR,
	TIEC440PVR,
	TIEC440USERRESET,
	TIEDCRBASEADDR,
	TRCC440TRACEDISABLE,
	TRCC440TRIGGEREVENTIN

);

parameter CLOCK_DELAY = "FALSE";
parameter DCR_AUTOLOCK_ENABLE = "TRUE";
parameter PPCDM_ASYNCMODE = "FALSE";
parameter PPCDS_ASYNCMODE = "FALSE";
parameter PPCS0_WIDTH_128N64 = "TRUE";
parameter PPCS1_WIDTH_128N64 = "TRUE";
parameter [0:16] APU_CONTROL = 17'h02000;
parameter [0:23] APU_UDI0 = 24'h000000;
parameter [0:23] APU_UDI1 = 24'h000000;
parameter [0:23] APU_UDI10 = 24'h000000;
parameter [0:23] APU_UDI11 = 24'h000000;
parameter [0:23] APU_UDI12 = 24'h000000;
parameter [0:23] APU_UDI13 = 24'h000000;
parameter [0:23] APU_UDI14 = 24'h000000;
parameter [0:23] APU_UDI15 = 24'h000000;
parameter [0:23] APU_UDI2 = 24'h000000;
parameter [0:23] APU_UDI3 = 24'h000000;
parameter [0:23] APU_UDI4 = 24'h000000;
parameter [0:23] APU_UDI5 = 24'h000000;
parameter [0:23] APU_UDI6 = 24'h000000;
parameter [0:23] APU_UDI7 = 24'h000000;
parameter [0:23] APU_UDI8 = 24'h000000;
parameter [0:23] APU_UDI9 = 24'h000000;
parameter [0:31] DMA0_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA0_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] INTERCONNECT_IMASK = 32'hFFFFFFFF;
parameter [0:31] INTERCONNECT_TMPL_SEL = 32'h3FFFFFFF;
parameter [0:31] MI_ARBCONFIG = 32'h00432010;
parameter [0:31] MI_BANKCONFLICT_MASK = 32'h00000000;
parameter [0:31] MI_CONTROL = 32'h0000008F;
parameter [0:31] MI_ROWCONFLICT_MASK = 32'h00000000;
parameter [0:31] PPCM_ARBCONFIG = 32'h00432010;
parameter [0:31] PPCM_CONTROL = 32'h8000009F;
parameter [0:31] PPCM_COUNTER = 32'h00000500;
parameter [0:31] PPCS0_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_CONTROL = 32'h8033336C;
parameter [0:31] PPCS1_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_CONTROL = 32'h8033336C;
parameter [0:31] XBAR_ADDRMAP_TMPL0 = 32'hFFFF0000;
parameter [0:31] XBAR_ADDRMAP_TMPL1 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL2 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL3 = 32'h00000000;
parameter [0:7] DMA0_CONTROL = 8'h00;
parameter [0:7] DMA1_CONTROL = 8'h00;
parameter [0:7] DMA2_CONTROL = 8'h00;
parameter [0:7] DMA3_CONTROL = 8'h00;
parameter [0:9] DMA0_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA0_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_TXIRQTIMER = 10'h3FF;

localparam in_delay = 1;
localparam out_delay = 0;
localparam CLK_DELAY = 0;

output APUFCMDECFPUOP;
output APUFCMDECLOAD;
output APUFCMDECNONAUTON;
output APUFCMDECSTORE;
output APUFCMDECUDIVALID;
output APUFCMENDIAN;
output APUFCMFLUSH;
output APUFCMINSTRVALID;
output APUFCMLOADDVALID;
output APUFCMMSRFE0;
output APUFCMMSRFE1;
output APUFCMNEXTINSTRREADY;
output APUFCMOPERANDVALID;
output APUFCMWRITEBACKOK;
output C440CPMCORESLEEPREQ;
output C440CPMDECIRPTREQ;
output C440CPMFITIRPTREQ;
output C440CPMMSRCE;
output C440CPMMSREE;
output C440CPMTIMERRESETREQ;
output C440CPMWDIRPTREQ;
output C440JTGTDO;
output C440JTGTDOEN;
output C440MACHINECHECK;
output C440RSTCHIPRESETREQ;
output C440RSTCORERESETREQ;
output C440RSTSYSTEMRESETREQ;
output C440TRCCYCLE;
output C440TRCTRIGGEREVENTOUT;
output DMA0LLRSTENGINEACK;
output DMA0LLRXDSTRDYN;
output DMA0LLTXEOFN;
output DMA0LLTXEOPN;
output DMA0LLTXSOFN;
output DMA0LLTXSOPN;
output DMA0LLTXSRCRDYN;
output DMA0RXIRQ;
output DMA0TXIRQ;
output DMA1LLRSTENGINEACK;
output DMA1LLRXDSTRDYN;
output DMA1LLTXEOFN;
output DMA1LLTXEOPN;
output DMA1LLTXSOFN;
output DMA1LLTXSOPN;
output DMA1LLTXSRCRDYN;
output DMA1RXIRQ;
output DMA1TXIRQ;
output DMA2LLRSTENGINEACK;
output DMA2LLRXDSTRDYN;
output DMA2LLTXEOFN;
output DMA2LLTXEOPN;
output DMA2LLTXSOFN;
output DMA2LLTXSOPN;
output DMA2LLTXSRCRDYN;
output DMA2RXIRQ;
output DMA2TXIRQ;
output DMA3LLRSTENGINEACK;
output DMA3LLRXDSTRDYN;
output DMA3LLTXEOFN;
output DMA3LLTXEOPN;
output DMA3LLTXSOFN;
output DMA3LLTXSOPN;
output DMA3LLTXSRCRDYN;
output DMA3RXIRQ;
output DMA3TXIRQ;
output MIMCADDRESSVALID;
output MIMCBANKCONFLICT;
output MIMCREADNOTWRITE;
output MIMCROWCONFLICT;
output MIMCWRITEDATAVALID;
output PPCCPMINTERCONNECTBUSY;
output PPCDMDCRREAD;
output PPCDMDCRWRITE;
output PPCDSDCRACK;
output PPCDSDCRTIMEOUTWAIT;
output PPCEICINTERCONNECTIRQ;
output PPCMPLBABORT;
output PPCMPLBBUSLOCK;
output PPCMPLBLOCKERR;
output PPCMPLBRDBURST;
output PPCMPLBREQUEST;
output PPCMPLBRNW;
output PPCMPLBWRBURST;
output PPCS0PLBADDRACK;
output PPCS0PLBRDBTERM;
output PPCS0PLBRDCOMP;
output PPCS0PLBRDDACK;
output PPCS0PLBREARBITRATE;
output PPCS0PLBWAIT;
output PPCS0PLBWRBTERM;
output PPCS0PLBWRCOMP;
output PPCS0PLBWRDACK;
output PPCS1PLBADDRACK;
output PPCS1PLBRDBTERM;
output PPCS1PLBRDCOMP;
output PPCS1PLBRDDACK;
output PPCS1PLBREARBITRATE;
output PPCS1PLBWAIT;
output PPCS1PLBWRBTERM;
output PPCS1PLBWRCOMP;
output PPCS1PLBWRDACK;
output [0:127] APUFCMLOADDATA;
output [0:127] MIMCWRITEDATA;
output [0:127] PPCMPLBWRDBUS;
output [0:127] PPCS0PLBRDDBUS;
output [0:127] PPCS1PLBRDDBUS;
output [0:13] C440TRCTRIGGEREVENTTYPE;
output [0:15] MIMCBYTEENABLE;
output [0:15] PPCMPLBBE;
output [0:15] PPCMPLBTATTRIBUTE;
output [0:1] PPCMPLBPRIORITY;
output [0:1] PPCS0PLBSSIZE;
output [0:1] PPCS1PLBSSIZE;
output [0:2] APUFCMDECLDSTXFERSIZE;
output [0:2] C440TRCBRANCHSTATUS;
output [0:2] PPCMPLBTYPE;
output [0:31] APUFCMINSTRUCTION;
output [0:31] APUFCMRADATA;
output [0:31] APUFCMRBDATA;
output [0:31] DMA0LLTXD;
output [0:31] DMA1LLTXD;
output [0:31] DMA2LLTXD;
output [0:31] DMA3LLTXD;
output [0:31] PPCDMDCRDBUSOUT;
output [0:31] PPCDSDCRDBUSIN;
output [0:31] PPCMPLBABUS;
output [0:35] MIMCADDRESS;
output [0:3] APUFCMDECUDI;
output [0:3] APUFCMLOADBYTEADDR;
output [0:3] DMA0LLTXREM;
output [0:3] DMA1LLTXREM;
output [0:3] DMA2LLTXREM;
output [0:3] DMA3LLTXREM;
output [0:3] PPCMPLBSIZE;
output [0:3] PPCS0PLBMBUSY;
output [0:3] PPCS0PLBMIRQ;
output [0:3] PPCS0PLBMRDERR;
output [0:3] PPCS0PLBMWRERR;
output [0:3] PPCS0PLBRDWDADDR;
output [0:3] PPCS1PLBMBUSY;
output [0:3] PPCS1PLBMIRQ;
output [0:3] PPCS1PLBMRDERR;
output [0:3] PPCS1PLBMWRERR;
output [0:3] PPCS1PLBRDWDADDR;
output [0:4] C440TRCEXECUTIONSTATUS;
output [0:6] C440TRCTRACESTATUS;
output [0:7] C440DBGSYSTEMCONTROL;
output [0:9] PPCDMDCRABUS;
output [20:21] PPCDMDCRUABUS;
output [28:31] PPCMPLBUABUS;

input CPMC440CLK;
input CPMC440CLKEN;
input CPMC440CORECLOCKINACTIVE;
input CPMC440TIMERCLOCK;
input CPMDCRCLK;
input CPMDMA0LLCLK;
input CPMDMA1LLCLK;
input CPMDMA2LLCLK;
input CPMDMA3LLCLK;
input CPMFCMCLK;
input CPMINTERCONNECTCLK;
input CPMINTERCONNECTCLKEN;
input CPMINTERCONNECTCLKNTO1;
input CPMMCCLK;
input CPMPPCMPLBCLK;
input CPMPPCS0PLBCLK;
input CPMPPCS1PLBCLK;
input DBGC440DEBUGHALT;
input DBGC440UNCONDDEBUGEVENT;
input DCRPPCDMACK;
input DCRPPCDMTIMEOUTWAIT;
input DCRPPCDSREAD;
input DCRPPCDSWRITE;
input EICC440CRITIRQ;
input EICC440EXTIRQ;
input FCMAPUCONFIRMINSTR;
input FCMAPUDONE;
input FCMAPUEXCEPTION;
input FCMAPUFPSCRFEX;
input FCMAPURESULTVALID;
input FCMAPUSLEEPNOTREADY;
input JTGC440TCK;
input JTGC440TDI;
input JTGC440TMS;
input JTGC440TRSTNEG;
input LLDMA0RSTENGINEREQ;
input LLDMA0RXEOFN;
input LLDMA0RXEOPN;
input LLDMA0RXSOFN;
input LLDMA0RXSOPN;
input LLDMA0RXSRCRDYN;
input LLDMA0TXDSTRDYN;
input LLDMA1RSTENGINEREQ;
input LLDMA1RXEOFN;
input LLDMA1RXEOPN;
input LLDMA1RXSOFN;
input LLDMA1RXSOPN;
input LLDMA1RXSRCRDYN;
input LLDMA1TXDSTRDYN;
input LLDMA2RSTENGINEREQ;
input LLDMA2RXEOFN;
input LLDMA2RXEOPN;
input LLDMA2RXSOFN;
input LLDMA2RXSOPN;
input LLDMA2RXSRCRDYN;
input LLDMA2TXDSTRDYN;
input LLDMA3RSTENGINEREQ;
input LLDMA3RXEOFN;
input LLDMA3RXEOPN;
input LLDMA3RXSOFN;
input LLDMA3RXSOPN;
input LLDMA3RXSRCRDYN;
input LLDMA3TXDSTRDYN;
input MCMIADDRREADYTOACCEPT;
input MCMIREADDATAERR;
input MCMIREADDATAVALID;
input PLBPPCMADDRACK;
input PLBPPCMMBUSY;
input PLBPPCMMIRQ;
input PLBPPCMMRDERR;
input PLBPPCMMWRERR;
input PLBPPCMRDBTERM;
input PLBPPCMRDDACK;
input PLBPPCMRDPENDREQ;
input PLBPPCMREARBITRATE;
input PLBPPCMTIMEOUT;
input PLBPPCMWRBTERM;
input PLBPPCMWRDACK;
input PLBPPCMWRPENDREQ;
input PLBPPCS0ABORT;
input PLBPPCS0BUSLOCK;
input PLBPPCS0LOCKERR;
input PLBPPCS0PAVALID;
input PLBPPCS0RDBURST;
input PLBPPCS0RDPENDREQ;
input PLBPPCS0RDPRIM;
input PLBPPCS0RNW;
input PLBPPCS0SAVALID;
input PLBPPCS0WRBURST;
input PLBPPCS0WRPENDREQ;
input PLBPPCS0WRPRIM;
input PLBPPCS1ABORT;
input PLBPPCS1BUSLOCK;
input PLBPPCS1LOCKERR;
input PLBPPCS1PAVALID;
input PLBPPCS1RDBURST;
input PLBPPCS1RDPENDREQ;
input PLBPPCS1RDPRIM;
input PLBPPCS1RNW;
input PLBPPCS1SAVALID;
input PLBPPCS1WRBURST;
input PLBPPCS1WRPENDREQ;
input PLBPPCS1WRPRIM;
input RSTC440RESETCHIP;
input RSTC440RESETCORE;
input RSTC440RESETSYSTEM;
input TIEC440ENDIANRESET;
input TRCC440TRACEDISABLE;
input TRCC440TRIGGEREVENTIN;
input [0:127] FCMAPUSTOREDATA;
input [0:127] MCMIREADDATA;
input [0:127] PLBPPCMRDDBUS;
input [0:127] PLBPPCS0WRDBUS;
input [0:127] PLBPPCS1WRDBUS;
input [0:15] PLBPPCS0BE;
input [0:15] PLBPPCS0TATTRIBUTE;
input [0:15] PLBPPCS1BE;
input [0:15] PLBPPCS1TATTRIBUTE;
input [0:1] PLBPPCMRDPENDPRI;
input [0:1] PLBPPCMREQPRI;
input [0:1] PLBPPCMSSIZE;
input [0:1] PLBPPCMWRPENDPRI;
input [0:1] PLBPPCS0MASTERID;
input [0:1] PLBPPCS0MSIZE;
input [0:1] PLBPPCS0RDPENDPRI;
input [0:1] PLBPPCS0REQPRI;
input [0:1] PLBPPCS0WRPENDPRI;
input [0:1] PLBPPCS1MASTERID;
input [0:1] PLBPPCS1MSIZE;
input [0:1] PLBPPCS1RDPENDPRI;
input [0:1] PLBPPCS1REQPRI;
input [0:1] PLBPPCS1WRPENDPRI;
input [0:1] TIEC440DCURDLDCACHEPLBPRIO;
input [0:1] TIEC440DCURDNONCACHEPLBPRIO;
input [0:1] TIEC440DCURDTOUCHPLBPRIO;
input [0:1] TIEC440DCURDURGENTPLBPRIO;
input [0:1] TIEC440DCUWRFLUSHPLBPRIO;
input [0:1] TIEC440DCUWRSTOREPLBPRIO;
input [0:1] TIEC440DCUWRURGENTPLBPRIO;
input [0:1] TIEC440ICURDFETCHPLBPRIO;
input [0:1] TIEC440ICURDSPECPLBPRIO;
input [0:1] TIEC440ICURDTOUCHPLBPRIO;
input [0:1] TIEDCRBASEADDR;
input [0:2] PLBPPCS0TYPE;
input [0:2] PLBPPCS1TYPE;
input [0:31] DCRPPCDMDBUSIN;
input [0:31] DCRPPCDSDBUSOUT;
input [0:31] FCMAPURESULT;
input [0:31] LLDMA0RXD;
input [0:31] LLDMA1RXD;
input [0:31] LLDMA2RXD;
input [0:31] LLDMA3RXD;
input [0:31] PLBPPCS0ABUS;
input [0:31] PLBPPCS1ABUS;
input [0:3] FCMAPUCR;
input [0:3] LLDMA0RXREM;
input [0:3] LLDMA1RXREM;
input [0:3] LLDMA2RXREM;
input [0:3] LLDMA3RXREM;
input [0:3] PLBPPCMRDWDADDR;
input [0:3] PLBPPCS0SIZE;
input [0:3] PLBPPCS1SIZE;
input [0:3] TIEC440ERPNRESET;
input [0:3] TIEC440USERRESET;
input [0:4] DBGC440SYSTEMSTATUS;
input [0:9] DCRPPCDSABUS;
input [28:31] PLBPPCS0UABUS;
input [28:31] PLBPPCS1UABUS;
input [28:31] TIEC440PIR;
input [28:31] TIEC440PVR;

reg [0:4] CLOCK_DELAY_BINARY;
reg DCR_AUTOLOCK_ENABLE_BINARY;
reg PPCDM_ASYNCMODE_BINARY;
reg PPCDS_ASYNCMODE_BINARY;
reg PPCS0_WIDTH_128N64_BINARY;
reg PPCS1_WIDTH_128N64_BINARY;

tri0 GSR = glbl.GSR;


initial begin
	case (PPCS0_WIDTH_128N64)
		"FALSE" : PPCS0_WIDTH_128N64_BINARY = 1'b0;
		"TRUE" : PPCS0_WIDTH_128N64_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCS0_WIDTH_128N64 on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCS0_WIDTH_128N64);
			$finish;
		end
	endcase

	case (PPCS1_WIDTH_128N64)
		"FALSE" : PPCS1_WIDTH_128N64_BINARY = 1'b0;
		"TRUE" : PPCS1_WIDTH_128N64_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCS1_WIDTH_128N64 on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCS1_WIDTH_128N64);
			$finish;
		end
	endcase

	case (PPCDM_ASYNCMODE)
		"FALSE" : PPCDM_ASYNCMODE_BINARY = 1'b0;
		"TRUE" : PPCDM_ASYNCMODE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCDM_ASYNCMODE on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCDM_ASYNCMODE);
			$finish;
		end
	endcase

	case (PPCDS_ASYNCMODE)
		"FALSE" : PPCDS_ASYNCMODE_BINARY = 1'b0;
		"TRUE" : PPCDS_ASYNCMODE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCDS_ASYNCMODE on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCDS_ASYNCMODE);
			$finish;
		end
	endcase

	case (DCR_AUTOLOCK_ENABLE)
		"FALSE" : DCR_AUTOLOCK_ENABLE_BINARY = 1'b0;
		"TRUE" : DCR_AUTOLOCK_ENABLE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute DCR_AUTOLOCK_ENABLE on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", DCR_AUTOLOCK_ENABLE);
			$finish;
		end
	endcase

	case (CLOCK_DELAY)
//		"FALSE" : CLOCK_DELAY_BINARY = 1'b0;
//		"TRUE" : CLOCK_DELAY_BINARY = 1'b1;
//		"FALSE" : CLOCK_DELAY_BINARY = 5'b00100;
		"FALSE" : CLOCK_DELAY_BINARY = 5'b10000;
		"TRUE" : CLOCK_DELAY_BINARY = 5'b00000;
		default : begin
			$display("Attribute Syntax Error : The Attribute CLOCK_DELAY on PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", CLOCK_DELAY);
			$finish;
		end
	endcase

end

wire APUFCMDECFPUOP_delay;
wire APUFCMDECLOAD_delay;
wire APUFCMDECNONAUTON_delay;
wire APUFCMDECSTORE_delay;
wire APUFCMDECUDIVALID_delay;
wire APUFCMENDIAN_delay;
wire APUFCMFLUSH_delay;
wire APUFCMINSTRVALID_delay;
wire APUFCMLOADDVALID_delay;
wire APUFCMMSRFE0_delay;
wire APUFCMMSRFE1_delay;
wire APUFCMNEXTINSTRREADY_delay;
wire APUFCMOPERANDVALID_delay;
wire APUFCMWRITEBACKOK_delay;
wire C440CPMCORESLEEPREQ_delay;
wire C440CPMDECIRPTREQ_delay;
wire C440CPMFITIRPTREQ_delay;
wire C440CPMMSRCE_delay;
wire C440CPMMSREE_delay;
wire C440CPMTIMERRESETREQ_delay;
wire C440CPMWDIRPTREQ_delay;
wire C440JTGTDOEN_delay;
wire C440JTGTDO_delay;
wire C440MACHINECHECK_delay;
wire C440RSTCHIPRESETREQ_delay;
wire C440RSTCORERESETREQ_delay;
wire C440RSTSYSTEMRESETREQ_delay;
wire C440TRCCYCLE_delay;
wire C440TRCTRIGGEREVENTOUT_delay;
wire DMA0LLRSTENGINEACK_delay;
wire DMA0LLRXDSTRDYN_delay;
wire DMA0LLTXEOFN_delay;
wire DMA0LLTXEOPN_delay;
wire DMA0LLTXSOFN_delay;
wire DMA0LLTXSOPN_delay;
wire DMA0LLTXSRCRDYN_delay;
wire DMA0RXIRQ_delay;
wire DMA0TXIRQ_delay;
wire DMA1LLRSTENGINEACK_delay;
wire DMA1LLRXDSTRDYN_delay;
wire DMA1LLTXEOFN_delay;
wire DMA1LLTXEOPN_delay;
wire DMA1LLTXSOFN_delay;
wire DMA1LLTXSOPN_delay;
wire DMA1LLTXSRCRDYN_delay;
wire DMA1RXIRQ_delay;
wire DMA1TXIRQ_delay;
wire DMA2LLRSTENGINEACK_delay;
wire DMA2LLRXDSTRDYN_delay;
wire DMA2LLTXEOFN_delay;
wire DMA2LLTXEOPN_delay;
wire DMA2LLTXSOFN_delay;
wire DMA2LLTXSOPN_delay;
wire DMA2LLTXSRCRDYN_delay;
wire DMA2RXIRQ_delay;
wire DMA2TXIRQ_delay;
wire DMA3LLRSTENGINEACK_delay;
wire DMA3LLRXDSTRDYN_delay;
wire DMA3LLTXEOFN_delay;
wire DMA3LLTXEOPN_delay;
wire DMA3LLTXSOFN_delay;
wire DMA3LLTXSOPN_delay;
wire DMA3LLTXSRCRDYN_delay;
wire DMA3RXIRQ_delay;
wire DMA3TXIRQ_delay;
wire MIMCADDRESSVALID_delay;
wire MIMCBANKCONFLICT_delay;
wire MIMCREADNOTWRITE_delay;
wire MIMCROWCONFLICT_delay;
wire MIMCWRITEDATAVALID_delay;
wire PPCCPMINTERCONNECTBUSY_delay;
wire PPCDMDCRREAD_delay;
wire PPCDMDCRWRITE_delay;
wire PPCDSDCRACK_delay;
wire PPCDSDCRTIMEOUTWAIT_delay;
wire PPCEICINTERCONNECTIRQ_delay;
wire PPCMPLBABORT_delay;
wire PPCMPLBBUSLOCK_delay;
wire PPCMPLBLOCKERR_delay;
wire PPCMPLBRDBURST_delay;
wire PPCMPLBREQUEST_delay;
wire PPCMPLBRNW_delay;
wire PPCMPLBWRBURST_delay;
wire PPCS0PLBADDRACK_delay;
wire PPCS0PLBRDBTERM_delay;
wire PPCS0PLBRDCOMP_delay;
wire PPCS0PLBRDDACK_delay;
wire PPCS0PLBREARBITRATE_delay;
wire PPCS0PLBWAIT_delay;
wire PPCS0PLBWRBTERM_delay;
wire PPCS0PLBWRCOMP_delay;
wire PPCS0PLBWRDACK_delay;
wire PPCS1PLBADDRACK_delay;
wire PPCS1PLBRDBTERM_delay;
wire PPCS1PLBRDCOMP_delay;
wire PPCS1PLBRDDACK_delay;
wire PPCS1PLBREARBITRATE_delay;
wire PPCS1PLBWAIT_delay;
wire PPCS1PLBWRBTERM_delay;
wire PPCS1PLBWRCOMP_delay;
wire PPCS1PLBWRDACK_delay;
wire [0:127] APUFCMLOADDATA_delay;
wire [0:127] MIMCWRITEDATA_delay;
wire [0:127] PPCMPLBWRDBUS_delay;
wire [0:127] PPCS0PLBRDDBUS_delay;
wire [0:127] PPCS1PLBRDDBUS_delay;
wire [0:13] C440TRCTRIGGEREVENTTYPE_delay;
wire [0:15] MIMCBYTEENABLE_delay;
wire [0:15] PPCMPLBBE_delay;
wire [0:15] PPCMPLBTATTRIBUTE_delay;
wire [0:1] PPCMPLBPRIORITY_delay;
wire [0:1] PPCS0PLBSSIZE_delay;
wire [0:1] PPCS1PLBSSIZE_delay;
wire [0:2] APUFCMDECLDSTXFERSIZE_delay;
wire [0:2] C440TRCBRANCHSTATUS_delay;
wire [0:2] PPCMPLBTYPE_delay;
wire [0:31] APUFCMINSTRUCTION_delay;
wire [0:31] APUFCMRADATA_delay;
wire [0:31] APUFCMRBDATA_delay;
wire [0:31] DMA0LLTXD_delay;
wire [0:31] DMA1LLTXD_delay;
wire [0:31] DMA2LLTXD_delay;
wire [0:31] DMA3LLTXD_delay;
wire [0:31] PPCDMDCRDBUSOUT_delay;
wire [0:31] PPCDSDCRDBUSIN_delay;
wire [0:31] PPCMPLBABUS_delay;
wire [0:35] MIMCADDRESS_delay;
wire [0:3] APUFCMDECUDI_delay;
wire [0:3] APUFCMLOADBYTEADDR_delay;
wire [0:3] DMA0LLTXREM_delay;
wire [0:3] DMA1LLTXREM_delay;
wire [0:3] DMA2LLTXREM_delay;
wire [0:3] DMA3LLTXREM_delay;
wire [0:3] PPCMPLBSIZE_delay;
wire [0:3] PPCS0PLBMBUSY_delay;
wire [0:3] PPCS0PLBMIRQ_delay;
wire [0:3] PPCS0PLBMRDERR_delay;
wire [0:3] PPCS0PLBMWRERR_delay;
wire [0:3] PPCS0PLBRDWDADDR_delay;
wire [0:3] PPCS1PLBMBUSY_delay;
wire [0:3] PPCS1PLBMIRQ_delay;
wire [0:3] PPCS1PLBMRDERR_delay;
wire [0:3] PPCS1PLBMWRERR_delay;
wire [0:3] PPCS1PLBRDWDADDR_delay;
wire [0:4] C440TRCEXECUTIONSTATUS_delay;
wire [0:6] C440TRCTRACESTATUS_delay;
wire [0:7] C440DBGSYSTEMCONTROL_delay;
wire [0:9] PPCDMDCRABUS_delay;
wire [20:21] PPCDMDCRUABUS_delay;
wire [28:31] PPCMPLBUABUS_delay;

wire CPMC440CLKEN_delay;
wire CPMC440CLK_delay;
wire CPMC440CORECLOCKINACTIVE_delay;
wire CPMC440TIMERCLOCK_delay;
wire CPMDCRCLK_delay;
wire CPMDMA0LLCLK_delay;
wire CPMDMA1LLCLK_delay;
wire CPMDMA2LLCLK_delay;
wire CPMDMA3LLCLK_delay;
wire CPMFCMCLK_delay;
wire CPMINTERCONNECTCLKEN_delay;
wire CPMINTERCONNECTCLKNTO1_delay;
wire CPMINTERCONNECTCLK_delay;
wire CPMMCCLK_delay;
wire CPMPPCMPLBCLK_delay;
wire CPMPPCS0PLBCLK_delay;
wire CPMPPCS1PLBCLK_delay;
wire DBGC440DEBUGHALT_delay;
wire DBGC440UNCONDDEBUGEVENT_delay;
wire DCRPPCDMACK_delay;
wire DCRPPCDMTIMEOUTWAIT_delay;
wire DCRPPCDSREAD_delay;
wire DCRPPCDSWRITE_delay;
wire EICC440CRITIRQ_delay;
wire EICC440EXTIRQ_delay;
wire FCMAPUCONFIRMINSTR_delay;
wire FCMAPUDONE_delay;
wire FCMAPUEXCEPTION_delay;
wire FCMAPUFPSCRFEX_delay;
wire FCMAPURESULTVALID_delay;
wire FCMAPUSLEEPNOTREADY_delay;
wire JTGC440TCK_delay;
wire JTGC440TDI_delay;
wire JTGC440TMS_delay;
wire JTGC440TRSTNEG_delay;
wire LLDMA0RSTENGINEREQ_delay;
wire LLDMA0RXEOFN_delay;
wire LLDMA0RXEOPN_delay;
wire LLDMA0RXSOFN_delay;
wire LLDMA0RXSOPN_delay;
wire LLDMA0RXSRCRDYN_delay;
wire LLDMA0TXDSTRDYN_delay;
wire LLDMA1RSTENGINEREQ_delay;
wire LLDMA1RXEOFN_delay;
wire LLDMA1RXEOPN_delay;
wire LLDMA1RXSOFN_delay;
wire LLDMA1RXSOPN_delay;
wire LLDMA1RXSRCRDYN_delay;
wire LLDMA1TXDSTRDYN_delay;
wire LLDMA2RSTENGINEREQ_delay;
wire LLDMA2RXEOFN_delay;
wire LLDMA2RXEOPN_delay;
wire LLDMA2RXSOFN_delay;
wire LLDMA2RXSOPN_delay;
wire LLDMA2RXSRCRDYN_delay;
wire LLDMA2TXDSTRDYN_delay;
wire LLDMA3RSTENGINEREQ_delay;
wire LLDMA3RXEOFN_delay;
wire LLDMA3RXEOPN_delay;
wire LLDMA3RXSOFN_delay;
wire LLDMA3RXSOPN_delay;
wire LLDMA3RXSRCRDYN_delay;
wire LLDMA3TXDSTRDYN_delay;
wire MCMIADDRREADYTOACCEPT_delay;
wire MCMIREADDATAERR_delay;
wire MCMIREADDATAVALID_delay;
wire PLBPPCMADDRACK_delay;
wire PLBPPCMMBUSY_delay;
wire PLBPPCMMIRQ_delay;
wire PLBPPCMMRDERR_delay;
wire PLBPPCMMWRERR_delay;
wire PLBPPCMRDBTERM_delay;
wire PLBPPCMRDDACK_delay;
wire PLBPPCMRDPENDREQ_delay;
wire PLBPPCMREARBITRATE_delay;
wire PLBPPCMTIMEOUT_delay;
wire PLBPPCMWRBTERM_delay;
wire PLBPPCMWRDACK_delay;
wire PLBPPCMWRPENDREQ_delay;
wire PLBPPCS0ABORT_delay;
wire PLBPPCS0BUSLOCK_delay;
wire PLBPPCS0LOCKERR_delay;
wire PLBPPCS0PAVALID_delay;
wire PLBPPCS0RDBURST_delay;
wire PLBPPCS0RDPENDREQ_delay;
wire PLBPPCS0RDPRIM_delay;
wire PLBPPCS0RNW_delay;
wire PLBPPCS0SAVALID_delay;
wire PLBPPCS0WRBURST_delay;
wire PLBPPCS0WRPENDREQ_delay;
wire PLBPPCS0WRPRIM_delay;
wire PLBPPCS1ABORT_delay;
wire PLBPPCS1BUSLOCK_delay;
wire PLBPPCS1LOCKERR_delay;
wire PLBPPCS1PAVALID_delay;
wire PLBPPCS1RDBURST_delay;
wire PLBPPCS1RDPENDREQ_delay;
wire PLBPPCS1RDPRIM_delay;
wire PLBPPCS1RNW_delay;
wire PLBPPCS1SAVALID_delay;
wire PLBPPCS1WRBURST_delay;
wire PLBPPCS1WRPENDREQ_delay;
wire PLBPPCS1WRPRIM_delay;
wire RSTC440RESETCHIP_delay;
wire RSTC440RESETCORE_delay;
wire RSTC440RESETSYSTEM_delay;
wire TIEC440ENDIANRESET_delay;
wire TRCC440TRACEDISABLE_delay;
wire TRCC440TRIGGEREVENTIN_delay;
wire [0:127] FCMAPUSTOREDATA_delay;
wire [0:127] MCMIREADDATA_delay;
wire [0:127] PLBPPCMRDDBUS_delay;
wire [0:127] PLBPPCS0WRDBUS_delay;
wire [0:127] PLBPPCS1WRDBUS_delay;
wire [0:15] PLBPPCS0BE_delay;
wire [0:15] PLBPPCS0TATTRIBUTE_delay;
wire [0:15] PLBPPCS1BE_delay;
wire [0:15] PLBPPCS1TATTRIBUTE_delay;
wire [0:1] PLBPPCMRDPENDPRI_delay;
wire [0:1] PLBPPCMREQPRI_delay;
wire [0:1] PLBPPCMSSIZE_delay;
wire [0:1] PLBPPCMWRPENDPRI_delay;
wire [0:1] PLBPPCS0MASTERID_delay;
wire [0:1] PLBPPCS0MSIZE_delay;
wire [0:1] PLBPPCS0RDPENDPRI_delay;
wire [0:1] PLBPPCS0REQPRI_delay;
wire [0:1] PLBPPCS0WRPENDPRI_delay;
wire [0:1] PLBPPCS1MASTERID_delay;
wire [0:1] PLBPPCS1MSIZE_delay;
wire [0:1] PLBPPCS1RDPENDPRI_delay;
wire [0:1] PLBPPCS1REQPRI_delay;
wire [0:1] PLBPPCS1WRPENDPRI_delay;
wire [0:1] TIEC440DCURDLDCACHEPLBPRIO_delay;
wire [0:1] TIEC440DCURDNONCACHEPLBPRIO_delay;
wire [0:1] TIEC440DCURDTOUCHPLBPRIO_delay;
wire [0:1] TIEC440DCURDURGENTPLBPRIO_delay;
wire [0:1] TIEC440DCUWRFLUSHPLBPRIO_delay;
wire [0:1] TIEC440DCUWRSTOREPLBPRIO_delay;
wire [0:1] TIEC440DCUWRURGENTPLBPRIO_delay;
wire [0:1] TIEC440ICURDFETCHPLBPRIO_delay;
wire [0:1] TIEC440ICURDSPECPLBPRIO_delay;
wire [0:1] TIEC440ICURDTOUCHPLBPRIO_delay;
wire [0:1] TIEDCRBASEADDR_delay;
wire [0:2] PLBPPCS0TYPE_delay;
wire [0:2] PLBPPCS1TYPE_delay;
wire [0:31] DCRPPCDMDBUSIN_delay;
wire [0:31] DCRPPCDSDBUSOUT_delay;
wire [0:31] FCMAPURESULT_delay;
wire [0:31] LLDMA0RXD_delay;
wire [0:31] LLDMA1RXD_delay;
wire [0:31] LLDMA2RXD_delay;
wire [0:31] LLDMA3RXD_delay;
wire [0:31] PLBPPCS0ABUS_delay;
wire [0:31] PLBPPCS1ABUS_delay;
wire [0:3] FCMAPUCR_delay;
wire [0:3] LLDMA0RXREM_delay;
wire [0:3] LLDMA1RXREM_delay;
wire [0:3] LLDMA2RXREM_delay;
wire [0:3] LLDMA3RXREM_delay;
wire [0:3] PLBPPCMRDWDADDR_delay;
wire [0:3] PLBPPCS0SIZE_delay;
wire [0:3] PLBPPCS1SIZE_delay;
wire [0:3] TIEC440ERPNRESET_delay;
wire [0:3] TIEC440USERRESET_delay;
wire [0:4] DBGC440SYSTEMSTATUS_delay;
wire [0:9] DCRPPCDSABUS_delay;
wire [28:31] PLBPPCS0UABUS_delay;
wire [28:31] PLBPPCS1UABUS_delay;
wire [28:31] TIEC440PIR_delay;
wire [28:31] TIEC440PVR_delay;


assign #(out_delay) APUFCMDECFPUOP = APUFCMDECFPUOP_delay;
assign #(out_delay) APUFCMDECLDSTXFERSIZE = APUFCMDECLDSTXFERSIZE_delay;
assign #(out_delay) APUFCMDECLOAD = APUFCMDECLOAD_delay;
assign #(out_delay) APUFCMDECNONAUTON = APUFCMDECNONAUTON_delay;
assign #(out_delay) APUFCMDECSTORE = APUFCMDECSTORE_delay;
assign #(out_delay) APUFCMDECUDI = APUFCMDECUDI_delay;
assign #(out_delay) APUFCMDECUDIVALID = APUFCMDECUDIVALID_delay;
assign #(out_delay) APUFCMENDIAN = APUFCMENDIAN_delay;
assign #(out_delay) APUFCMFLUSH = APUFCMFLUSH_delay;
assign #(out_delay) APUFCMINSTRUCTION = APUFCMINSTRUCTION_delay;
assign #(out_delay) APUFCMINSTRVALID = APUFCMINSTRVALID_delay;
assign #(out_delay) APUFCMLOADBYTEADDR = APUFCMLOADBYTEADDR_delay;
assign #(out_delay) APUFCMLOADDATA = APUFCMLOADDATA_delay;
assign #(out_delay) APUFCMLOADDVALID = APUFCMLOADDVALID_delay;
assign #(out_delay) APUFCMMSRFE0 = APUFCMMSRFE0_delay;
assign #(out_delay) APUFCMMSRFE1 = APUFCMMSRFE1_delay;
assign #(out_delay) APUFCMNEXTINSTRREADY = APUFCMNEXTINSTRREADY_delay;
assign #(out_delay) APUFCMOPERANDVALID = APUFCMOPERANDVALID_delay;
assign #(out_delay) APUFCMRADATA = APUFCMRADATA_delay;
assign #(out_delay) APUFCMRBDATA = APUFCMRBDATA_delay;
assign #(out_delay) APUFCMWRITEBACKOK = APUFCMWRITEBACKOK_delay;
assign #(out_delay) C440CPMCORESLEEPREQ = C440CPMCORESLEEPREQ_delay;
assign #(out_delay) C440CPMDECIRPTREQ = C440CPMDECIRPTREQ_delay;
assign #(out_delay) C440CPMFITIRPTREQ = C440CPMFITIRPTREQ_delay;
assign #(out_delay) C440CPMMSRCE = C440CPMMSRCE_delay;
assign #(out_delay) C440CPMMSREE = C440CPMMSREE_delay;
assign #(out_delay) C440CPMTIMERRESETREQ = C440CPMTIMERRESETREQ_delay;
assign #(out_delay) C440CPMWDIRPTREQ = C440CPMWDIRPTREQ_delay;
assign #(out_delay) C440DBGSYSTEMCONTROL = C440DBGSYSTEMCONTROL_delay;
assign #(out_delay) C440JTGTDO = C440JTGTDO_delay;
assign #(out_delay) C440JTGTDOEN = C440JTGTDOEN_delay;
assign #(out_delay) C440MACHINECHECK = C440MACHINECHECK_delay;
assign #(out_delay) C440RSTCHIPRESETREQ = C440RSTCHIPRESETREQ_delay;
assign #(out_delay) C440RSTCORERESETREQ = C440RSTCORERESETREQ_delay;
assign #(out_delay) C440RSTSYSTEMRESETREQ = C440RSTSYSTEMRESETREQ_delay;
assign #(out_delay) C440TRCBRANCHSTATUS = C440TRCBRANCHSTATUS_delay;
assign #(out_delay) C440TRCCYCLE = C440TRCCYCLE_delay;
assign #(out_delay) C440TRCEXECUTIONSTATUS = C440TRCEXECUTIONSTATUS_delay;
assign #(out_delay) C440TRCTRACESTATUS = C440TRCTRACESTATUS_delay;
assign #(out_delay) C440TRCTRIGGEREVENTOUT = C440TRCTRIGGEREVENTOUT_delay;
assign #(out_delay) C440TRCTRIGGEREVENTTYPE = C440TRCTRIGGEREVENTTYPE_delay;
assign #(out_delay) DMA0LLRSTENGINEACK = DMA0LLRSTENGINEACK_delay;
assign #(out_delay) DMA0LLRXDSTRDYN = DMA0LLRXDSTRDYN_delay;
assign #(out_delay) DMA0LLTXD = DMA0LLTXD_delay;
assign #(out_delay) DMA0LLTXEOFN = DMA0LLTXEOFN_delay;
assign #(out_delay) DMA0LLTXEOPN = DMA0LLTXEOPN_delay;
assign #(out_delay) DMA0LLTXREM = DMA0LLTXREM_delay;
assign #(out_delay) DMA0LLTXSOFN = DMA0LLTXSOFN_delay;
assign #(out_delay) DMA0LLTXSOPN = DMA0LLTXSOPN_delay;
assign #(out_delay) DMA0LLTXSRCRDYN = DMA0LLTXSRCRDYN_delay;
assign #(out_delay) DMA0RXIRQ = DMA0RXIRQ_delay;
assign #(out_delay) DMA0TXIRQ = DMA0TXIRQ_delay;
assign #(out_delay) DMA1LLRSTENGINEACK = DMA1LLRSTENGINEACK_delay;
assign #(out_delay) DMA1LLRXDSTRDYN = DMA1LLRXDSTRDYN_delay;
assign #(out_delay) DMA1LLTXD = DMA1LLTXD_delay;
assign #(out_delay) DMA1LLTXEOFN = DMA1LLTXEOFN_delay;
assign #(out_delay) DMA1LLTXEOPN = DMA1LLTXEOPN_delay;
assign #(out_delay) DMA1LLTXREM = DMA1LLTXREM_delay;
assign #(out_delay) DMA1LLTXSOFN = DMA1LLTXSOFN_delay;
assign #(out_delay) DMA1LLTXSOPN = DMA1LLTXSOPN_delay;
assign #(out_delay) DMA1LLTXSRCRDYN = DMA1LLTXSRCRDYN_delay;
assign #(out_delay) DMA1RXIRQ = DMA1RXIRQ_delay;
assign #(out_delay) DMA1TXIRQ = DMA1TXIRQ_delay;
assign #(out_delay) DMA2LLRSTENGINEACK = DMA2LLRSTENGINEACK_delay;
assign #(out_delay) DMA2LLRXDSTRDYN = DMA2LLRXDSTRDYN_delay;
assign #(out_delay) DMA2LLTXD = DMA2LLTXD_delay;
assign #(out_delay) DMA2LLTXEOFN = DMA2LLTXEOFN_delay;
assign #(out_delay) DMA2LLTXEOPN = DMA2LLTXEOPN_delay;
assign #(out_delay) DMA2LLTXREM = DMA2LLTXREM_delay;
assign #(out_delay) DMA2LLTXSOFN = DMA2LLTXSOFN_delay;
assign #(out_delay) DMA2LLTXSOPN = DMA2LLTXSOPN_delay;
assign #(out_delay) DMA2LLTXSRCRDYN = DMA2LLTXSRCRDYN_delay;
assign #(out_delay) DMA2RXIRQ = DMA2RXIRQ_delay;
assign #(out_delay) DMA2TXIRQ = DMA2TXIRQ_delay;
assign #(out_delay) DMA3LLRSTENGINEACK = DMA3LLRSTENGINEACK_delay;
assign #(out_delay) DMA3LLRXDSTRDYN = DMA3LLRXDSTRDYN_delay;
assign #(out_delay) DMA3LLTXD = DMA3LLTXD_delay;
assign #(out_delay) DMA3LLTXEOFN = DMA3LLTXEOFN_delay;
assign #(out_delay) DMA3LLTXEOPN = DMA3LLTXEOPN_delay;
assign #(out_delay) DMA3LLTXREM = DMA3LLTXREM_delay;
assign #(out_delay) DMA3LLTXSOFN = DMA3LLTXSOFN_delay;
assign #(out_delay) DMA3LLTXSOPN = DMA3LLTXSOPN_delay;
assign #(out_delay) DMA3LLTXSRCRDYN = DMA3LLTXSRCRDYN_delay;
assign #(out_delay) DMA3RXIRQ = DMA3RXIRQ_delay;
assign #(out_delay) DMA3TXIRQ = DMA3TXIRQ_delay;
assign #(out_delay) MIMCADDRESS = MIMCADDRESS_delay;
assign #(out_delay) MIMCADDRESSVALID = MIMCADDRESSVALID_delay;
assign #(out_delay) MIMCBANKCONFLICT = MIMCBANKCONFLICT_delay;
assign #(out_delay) MIMCBYTEENABLE = MIMCBYTEENABLE_delay;
assign #(out_delay) MIMCREADNOTWRITE = MIMCREADNOTWRITE_delay;
assign #(out_delay) MIMCROWCONFLICT = MIMCROWCONFLICT_delay;
assign #(out_delay) MIMCWRITEDATA = MIMCWRITEDATA_delay;
assign #(out_delay) MIMCWRITEDATAVALID = MIMCWRITEDATAVALID_delay;
assign #(out_delay) PPCCPMINTERCONNECTBUSY = PPCCPMINTERCONNECTBUSY_delay;
assign #(out_delay) PPCDMDCRABUS = PPCDMDCRABUS_delay;
assign #(out_delay) PPCDMDCRDBUSOUT = PPCDMDCRDBUSOUT_delay;
assign #(out_delay) PPCDMDCRREAD = PPCDMDCRREAD_delay;
assign #(out_delay) PPCDMDCRUABUS = PPCDMDCRUABUS_delay;
assign #(out_delay) PPCDMDCRWRITE = PPCDMDCRWRITE_delay;
assign #(out_delay) PPCDSDCRACK = PPCDSDCRACK_delay;
assign #(out_delay) PPCDSDCRDBUSIN = PPCDSDCRDBUSIN_delay;
assign #(out_delay) PPCDSDCRTIMEOUTWAIT = PPCDSDCRTIMEOUTWAIT_delay;
assign #(out_delay) PPCEICINTERCONNECTIRQ = PPCEICINTERCONNECTIRQ_delay;
assign #(out_delay) PPCMPLBABORT = PPCMPLBABORT_delay;
assign #(out_delay) PPCMPLBABUS = PPCMPLBABUS_delay;
assign #(out_delay) PPCMPLBBE = PPCMPLBBE_delay;
assign #(out_delay) PPCMPLBBUSLOCK = PPCMPLBBUSLOCK_delay;
assign #(out_delay) PPCMPLBLOCKERR = PPCMPLBLOCKERR_delay;
assign #(out_delay) PPCMPLBPRIORITY = PPCMPLBPRIORITY_delay;
assign #(out_delay) PPCMPLBRDBURST = PPCMPLBRDBURST_delay;
assign #(out_delay) PPCMPLBREQUEST = PPCMPLBREQUEST_delay;
assign #(out_delay) PPCMPLBRNW = PPCMPLBRNW_delay;
assign #(out_delay) PPCMPLBSIZE = PPCMPLBSIZE_delay;
assign #(out_delay) PPCMPLBTATTRIBUTE = PPCMPLBTATTRIBUTE_delay;
assign #(out_delay) PPCMPLBTYPE = PPCMPLBTYPE_delay;
assign #(out_delay) PPCMPLBUABUS = PPCMPLBUABUS_delay;
assign #(out_delay) PPCMPLBWRBURST = PPCMPLBWRBURST_delay;
assign #(out_delay) PPCMPLBWRDBUS = PPCMPLBWRDBUS_delay;
assign #(out_delay) PPCS0PLBADDRACK = PPCS0PLBADDRACK_delay;
assign #(out_delay) PPCS0PLBMBUSY = PPCS0PLBMBUSY_delay;
assign #(out_delay) PPCS0PLBMIRQ = PPCS0PLBMIRQ_delay;
assign #(out_delay) PPCS0PLBMRDERR = PPCS0PLBMRDERR_delay;
assign #(out_delay) PPCS0PLBMWRERR = PPCS0PLBMWRERR_delay;
assign #(out_delay) PPCS0PLBRDBTERM = PPCS0PLBRDBTERM_delay;
assign #(out_delay) PPCS0PLBRDCOMP = PPCS0PLBRDCOMP_delay;
assign #(out_delay) PPCS0PLBRDDACK = PPCS0PLBRDDACK_delay;
assign #(out_delay) PPCS0PLBRDDBUS = PPCS0PLBRDDBUS_delay;
assign #(out_delay) PPCS0PLBRDWDADDR = PPCS0PLBRDWDADDR_delay;
assign #(out_delay) PPCS0PLBREARBITRATE = PPCS0PLBREARBITRATE_delay;
assign #(out_delay) PPCS0PLBSSIZE = PPCS0PLBSSIZE_delay;
assign #(out_delay) PPCS0PLBWAIT = PPCS0PLBWAIT_delay;
assign #(out_delay) PPCS0PLBWRBTERM = PPCS0PLBWRBTERM_delay;
assign #(out_delay) PPCS0PLBWRCOMP = PPCS0PLBWRCOMP_delay;
assign #(out_delay) PPCS0PLBWRDACK = PPCS0PLBWRDACK_delay;
assign #(out_delay) PPCS1PLBADDRACK = PPCS1PLBADDRACK_delay;
assign #(out_delay) PPCS1PLBMBUSY = PPCS1PLBMBUSY_delay;
assign #(out_delay) PPCS1PLBMIRQ = PPCS1PLBMIRQ_delay;
assign #(out_delay) PPCS1PLBMRDERR = PPCS1PLBMRDERR_delay;
assign #(out_delay) PPCS1PLBMWRERR = PPCS1PLBMWRERR_delay;
assign #(out_delay) PPCS1PLBRDBTERM = PPCS1PLBRDBTERM_delay;
assign #(out_delay) PPCS1PLBRDCOMP = PPCS1PLBRDCOMP_delay;
assign #(out_delay) PPCS1PLBRDDACK = PPCS1PLBRDDACK_delay;
assign #(out_delay) PPCS1PLBRDDBUS = PPCS1PLBRDDBUS_delay;
assign #(out_delay) PPCS1PLBRDWDADDR = PPCS1PLBRDWDADDR_delay;
assign #(out_delay) PPCS1PLBREARBITRATE = PPCS1PLBREARBITRATE_delay;
assign #(out_delay) PPCS1PLBSSIZE = PPCS1PLBSSIZE_delay;
assign #(out_delay) PPCS1PLBWAIT = PPCS1PLBWAIT_delay;
assign #(out_delay) PPCS1PLBWRBTERM = PPCS1PLBWRBTERM_delay;
assign #(out_delay) PPCS1PLBWRCOMP = PPCS1PLBWRCOMP_delay;
assign #(out_delay) PPCS1PLBWRDACK = PPCS1PLBWRDACK_delay;

assign #(CLK_DELAY) CPMC440CLK_delay = CPMC440CLK;
assign #(CLK_DELAY) CPMC440TIMERCLOCK_delay = CPMC440TIMERCLOCK;
assign #(CLK_DELAY) CPMDCRCLK_delay = CPMDCRCLK;
assign #(CLK_DELAY) CPMDMA0LLCLK_delay = CPMDMA0LLCLK;
assign #(CLK_DELAY) CPMDMA1LLCLK_delay = CPMDMA1LLCLK;
assign #(CLK_DELAY) CPMDMA2LLCLK_delay = CPMDMA2LLCLK;
assign #(CLK_DELAY) CPMDMA3LLCLK_delay = CPMDMA3LLCLK;
assign #(CLK_DELAY) CPMFCMCLK_delay = CPMFCMCLK;
assign #(CLK_DELAY) CPMINTERCONNECTCLK_delay = CPMINTERCONNECTCLK;
assign #(CLK_DELAY) CPMMCCLK_delay = CPMMCCLK;
assign #(CLK_DELAY) CPMPPCMPLBCLK_delay = CPMPPCMPLBCLK;
assign #(CLK_DELAY) CPMPPCS0PLBCLK_delay = CPMPPCS0PLBCLK;
assign #(CLK_DELAY) CPMPPCS1PLBCLK_delay = CPMPPCS1PLBCLK;
assign #(CLK_DELAY) JTGC440TCK_delay = JTGC440TCK;

assign #(in_delay) CPMC440CLKEN_delay = CPMC440CLKEN;
assign #(in_delay) CPMC440CORECLOCKINACTIVE_delay = CPMC440CORECLOCKINACTIVE;
assign #(in_delay) CPMINTERCONNECTCLKEN_delay = CPMINTERCONNECTCLKEN;
assign #(in_delay) CPMINTERCONNECTCLKNTO1_delay = CPMINTERCONNECTCLKNTO1;
assign #(in_delay) DBGC440DEBUGHALT_delay = DBGC440DEBUGHALT;
assign #(in_delay) DBGC440SYSTEMSTATUS_delay = DBGC440SYSTEMSTATUS;
assign #(in_delay) DBGC440UNCONDDEBUGEVENT_delay = DBGC440UNCONDDEBUGEVENT;
assign #(in_delay) DCRPPCDMACK_delay = DCRPPCDMACK;
assign #(in_delay) DCRPPCDMDBUSIN_delay = DCRPPCDMDBUSIN;
assign #(in_delay) DCRPPCDMTIMEOUTWAIT_delay = DCRPPCDMTIMEOUTWAIT;
assign #(in_delay) DCRPPCDSABUS_delay = DCRPPCDSABUS;
assign #(in_delay) DCRPPCDSDBUSOUT_delay = DCRPPCDSDBUSOUT;
assign #(in_delay) DCRPPCDSREAD_delay = DCRPPCDSREAD;
assign #(in_delay) DCRPPCDSWRITE_delay = DCRPPCDSWRITE;
assign #(in_delay) EICC440CRITIRQ_delay = EICC440CRITIRQ;
assign #(in_delay) EICC440EXTIRQ_delay = EICC440EXTIRQ;
assign #(in_delay) FCMAPUCONFIRMINSTR_delay = FCMAPUCONFIRMINSTR;
assign #(in_delay) FCMAPUCR_delay = FCMAPUCR;
assign #(in_delay) FCMAPUDONE_delay = FCMAPUDONE;
assign #(in_delay) FCMAPUEXCEPTION_delay = FCMAPUEXCEPTION;
assign #(in_delay) FCMAPUFPSCRFEX_delay = FCMAPUFPSCRFEX;
assign #(in_delay) FCMAPURESULTVALID_delay = FCMAPURESULTVALID;
assign #(in_delay) FCMAPURESULT_delay = FCMAPURESULT;
assign #(in_delay) FCMAPUSLEEPNOTREADY_delay = FCMAPUSLEEPNOTREADY;
assign #(in_delay) FCMAPUSTOREDATA_delay = FCMAPUSTOREDATA;
assign #(in_delay) JTGC440TDI_delay = JTGC440TDI;
assign #(in_delay) JTGC440TMS_delay = JTGC440TMS;
assign #(in_delay) JTGC440TRSTNEG_delay = JTGC440TRSTNEG;
assign #(in_delay) LLDMA0RSTENGINEREQ_delay = LLDMA0RSTENGINEREQ;
assign #(in_delay) LLDMA0RXD_delay = LLDMA0RXD;
assign #(in_delay) LLDMA0RXEOFN_delay = LLDMA0RXEOFN;
assign #(in_delay) LLDMA0RXEOPN_delay = LLDMA0RXEOPN;
assign #(in_delay) LLDMA0RXREM_delay = LLDMA0RXREM;
assign #(in_delay) LLDMA0RXSOFN_delay = LLDMA0RXSOFN;
assign #(in_delay) LLDMA0RXSOPN_delay = LLDMA0RXSOPN;
assign #(in_delay) LLDMA0RXSRCRDYN_delay = LLDMA0RXSRCRDYN;
assign #(in_delay) LLDMA0TXDSTRDYN_delay = LLDMA0TXDSTRDYN;
assign #(in_delay) LLDMA1RSTENGINEREQ_delay = LLDMA1RSTENGINEREQ;
assign #(in_delay) LLDMA1RXD_delay = LLDMA1RXD;
assign #(in_delay) LLDMA1RXEOFN_delay = LLDMA1RXEOFN;
assign #(in_delay) LLDMA1RXEOPN_delay = LLDMA1RXEOPN;
assign #(in_delay) LLDMA1RXREM_delay = LLDMA1RXREM;
assign #(in_delay) LLDMA1RXSOFN_delay = LLDMA1RXSOFN;
assign #(in_delay) LLDMA1RXSOPN_delay = LLDMA1RXSOPN;
assign #(in_delay) LLDMA1RXSRCRDYN_delay = LLDMA1RXSRCRDYN;
assign #(in_delay) LLDMA1TXDSTRDYN_delay = LLDMA1TXDSTRDYN;
assign #(in_delay) LLDMA2RSTENGINEREQ_delay = LLDMA2RSTENGINEREQ;
assign #(in_delay) LLDMA2RXD_delay = LLDMA2RXD;
assign #(in_delay) LLDMA2RXEOFN_delay = LLDMA2RXEOFN;
assign #(in_delay) LLDMA2RXEOPN_delay = LLDMA2RXEOPN;
assign #(in_delay) LLDMA2RXREM_delay = LLDMA2RXREM;
assign #(in_delay) LLDMA2RXSOFN_delay = LLDMA2RXSOFN;
assign #(in_delay) LLDMA2RXSOPN_delay = LLDMA2RXSOPN;
assign #(in_delay) LLDMA2RXSRCRDYN_delay = LLDMA2RXSRCRDYN;
assign #(in_delay) LLDMA2TXDSTRDYN_delay = LLDMA2TXDSTRDYN;
assign #(in_delay) LLDMA3RSTENGINEREQ_delay = LLDMA3RSTENGINEREQ;
assign #(in_delay) LLDMA3RXD_delay = LLDMA3RXD;
assign #(in_delay) LLDMA3RXEOFN_delay = LLDMA3RXEOFN;
assign #(in_delay) LLDMA3RXEOPN_delay = LLDMA3RXEOPN;
assign #(in_delay) LLDMA3RXREM_delay = LLDMA3RXREM;
assign #(in_delay) LLDMA3RXSOFN_delay = LLDMA3RXSOFN;
assign #(in_delay) LLDMA3RXSOPN_delay = LLDMA3RXSOPN;
assign #(in_delay) LLDMA3RXSRCRDYN_delay = LLDMA3RXSRCRDYN;
assign #(in_delay) LLDMA3TXDSTRDYN_delay = LLDMA3TXDSTRDYN;
assign #(in_delay) MCMIADDRREADYTOACCEPT_delay = MCMIADDRREADYTOACCEPT;
assign #(in_delay) MCMIREADDATAERR_delay = MCMIREADDATAERR;
assign #(in_delay) MCMIREADDATAVALID_delay = MCMIREADDATAVALID;
assign #(in_delay) MCMIREADDATA_delay = MCMIREADDATA;
assign #(in_delay) PLBPPCMADDRACK_delay = PLBPPCMADDRACK;
assign #(in_delay) PLBPPCMMBUSY_delay = PLBPPCMMBUSY;
assign #(in_delay) PLBPPCMMIRQ_delay = PLBPPCMMIRQ;
assign #(in_delay) PLBPPCMMRDERR_delay = PLBPPCMMRDERR;
assign #(in_delay) PLBPPCMMWRERR_delay = PLBPPCMMWRERR;
assign #(in_delay) PLBPPCMRDBTERM_delay = PLBPPCMRDBTERM;
assign #(in_delay) PLBPPCMRDDACK_delay = PLBPPCMRDDACK;
assign #(in_delay) PLBPPCMRDDBUS_delay = PLBPPCMRDDBUS;
assign #(in_delay) PLBPPCMRDPENDPRI_delay = PLBPPCMRDPENDPRI;
assign #(in_delay) PLBPPCMRDPENDREQ_delay = PLBPPCMRDPENDREQ;
assign #(in_delay) PLBPPCMRDWDADDR_delay = PLBPPCMRDWDADDR;
assign #(in_delay) PLBPPCMREARBITRATE_delay = PLBPPCMREARBITRATE;
assign #(in_delay) PLBPPCMREQPRI_delay = PLBPPCMREQPRI;
assign #(in_delay) PLBPPCMSSIZE_delay = PLBPPCMSSIZE;
assign #(in_delay) PLBPPCMTIMEOUT_delay = PLBPPCMTIMEOUT;
assign #(in_delay) PLBPPCMWRBTERM_delay = PLBPPCMWRBTERM;
assign #(in_delay) PLBPPCMWRDACK_delay = PLBPPCMWRDACK;
assign #(in_delay) PLBPPCMWRPENDPRI_delay = PLBPPCMWRPENDPRI;
assign #(in_delay) PLBPPCMWRPENDREQ_delay = PLBPPCMWRPENDREQ;
assign #(in_delay) PLBPPCS0ABORT_delay = PLBPPCS0ABORT;
assign #(in_delay) PLBPPCS0ABUS_delay = PLBPPCS0ABUS;
assign #(in_delay) PLBPPCS0BE_delay = PLBPPCS0BE;
assign #(in_delay) PLBPPCS0BUSLOCK_delay = PLBPPCS0BUSLOCK;
assign #(in_delay) PLBPPCS0LOCKERR_delay = PLBPPCS0LOCKERR;
assign #(in_delay) PLBPPCS0MASTERID_delay = PLBPPCS0MASTERID;
assign #(in_delay) PLBPPCS0MSIZE_delay = PLBPPCS0MSIZE;
assign #(in_delay) PLBPPCS0PAVALID_delay = PLBPPCS0PAVALID;
assign #(in_delay) PLBPPCS0RDBURST_delay = PLBPPCS0RDBURST;
assign #(in_delay) PLBPPCS0RDPENDPRI_delay = PLBPPCS0RDPENDPRI;
assign #(in_delay) PLBPPCS0RDPENDREQ_delay = PLBPPCS0RDPENDREQ;
assign #(in_delay) PLBPPCS0RDPRIM_delay = PLBPPCS0RDPRIM;
assign #(in_delay) PLBPPCS0REQPRI_delay = PLBPPCS0REQPRI;
assign #(in_delay) PLBPPCS0RNW_delay = PLBPPCS0RNW;
assign #(in_delay) PLBPPCS0SAVALID_delay = PLBPPCS0SAVALID;
assign #(in_delay) PLBPPCS0SIZE_delay = PLBPPCS0SIZE;
assign #(in_delay) PLBPPCS0TATTRIBUTE_delay = PLBPPCS0TATTRIBUTE;
assign #(in_delay) PLBPPCS0TYPE_delay = PLBPPCS0TYPE;
assign #(in_delay) PLBPPCS0UABUS_delay = PLBPPCS0UABUS;
assign #(in_delay) PLBPPCS0WRBURST_delay = PLBPPCS0WRBURST;
assign #(in_delay) PLBPPCS0WRDBUS_delay = PLBPPCS0WRDBUS;
assign #(in_delay) PLBPPCS0WRPENDPRI_delay = PLBPPCS0WRPENDPRI;
assign #(in_delay) PLBPPCS0WRPENDREQ_delay = PLBPPCS0WRPENDREQ;
assign #(in_delay) PLBPPCS0WRPRIM_delay = PLBPPCS0WRPRIM;
assign #(in_delay) PLBPPCS1ABORT_delay = PLBPPCS1ABORT;
assign #(in_delay) PLBPPCS1ABUS_delay = PLBPPCS1ABUS;
assign #(in_delay) PLBPPCS1BE_delay = PLBPPCS1BE;
assign #(in_delay) PLBPPCS1BUSLOCK_delay = PLBPPCS1BUSLOCK;
assign #(in_delay) PLBPPCS1LOCKERR_delay = PLBPPCS1LOCKERR;
assign #(in_delay) PLBPPCS1MASTERID_delay = PLBPPCS1MASTERID;
assign #(in_delay) PLBPPCS1MSIZE_delay = PLBPPCS1MSIZE;
assign #(in_delay) PLBPPCS1PAVALID_delay = PLBPPCS1PAVALID;
assign #(in_delay) PLBPPCS1RDBURST_delay = PLBPPCS1RDBURST;
assign #(in_delay) PLBPPCS1RDPENDPRI_delay = PLBPPCS1RDPENDPRI;
assign #(in_delay) PLBPPCS1RDPENDREQ_delay = PLBPPCS1RDPENDREQ;
assign #(in_delay) PLBPPCS1RDPRIM_delay = PLBPPCS1RDPRIM;
assign #(in_delay) PLBPPCS1REQPRI_delay = PLBPPCS1REQPRI;
assign #(in_delay) PLBPPCS1RNW_delay = PLBPPCS1RNW;
assign #(in_delay) PLBPPCS1SAVALID_delay = PLBPPCS1SAVALID;
assign #(in_delay) PLBPPCS1SIZE_delay = PLBPPCS1SIZE;
assign #(in_delay) PLBPPCS1TATTRIBUTE_delay = PLBPPCS1TATTRIBUTE;
assign #(in_delay) PLBPPCS1TYPE_delay = PLBPPCS1TYPE;
assign #(in_delay) PLBPPCS1UABUS_delay = PLBPPCS1UABUS;
assign #(in_delay) PLBPPCS1WRBURST_delay = PLBPPCS1WRBURST;
assign #(in_delay) PLBPPCS1WRDBUS_delay = PLBPPCS1WRDBUS;
assign #(in_delay) PLBPPCS1WRPENDPRI_delay = PLBPPCS1WRPENDPRI;
assign #(in_delay) PLBPPCS1WRPENDREQ_delay = PLBPPCS1WRPENDREQ;
assign #(in_delay) PLBPPCS1WRPRIM_delay = PLBPPCS1WRPRIM;
assign #(in_delay) RSTC440RESETCHIP_delay = RSTC440RESETCHIP;
assign #(in_delay) RSTC440RESETCORE_delay = RSTC440RESETCORE;
assign #(in_delay) RSTC440RESETSYSTEM_delay = RSTC440RESETSYSTEM;
assign #(in_delay) TIEC440DCURDLDCACHEPLBPRIO_delay = TIEC440DCURDLDCACHEPLBPRIO;
assign #(in_delay) TIEC440DCURDNONCACHEPLBPRIO_delay = TIEC440DCURDNONCACHEPLBPRIO;
assign #(in_delay) TIEC440DCURDTOUCHPLBPRIO_delay = TIEC440DCURDTOUCHPLBPRIO;
assign #(in_delay) TIEC440DCURDURGENTPLBPRIO_delay = TIEC440DCURDURGENTPLBPRIO;
assign #(in_delay) TIEC440DCUWRFLUSHPLBPRIO_delay = TIEC440DCUWRFLUSHPLBPRIO;
assign #(in_delay) TIEC440DCUWRSTOREPLBPRIO_delay = TIEC440DCUWRSTOREPLBPRIO;
assign #(in_delay) TIEC440DCUWRURGENTPLBPRIO_delay = TIEC440DCUWRURGENTPLBPRIO;
assign #(in_delay) TIEC440ENDIANRESET_delay = TIEC440ENDIANRESET;
assign #(in_delay) TIEC440ERPNRESET_delay = TIEC440ERPNRESET;
assign #(in_delay) TIEC440ICURDFETCHPLBPRIO_delay = TIEC440ICURDFETCHPLBPRIO;
assign #(in_delay) TIEC440ICURDSPECPLBPRIO_delay = TIEC440ICURDSPECPLBPRIO;
assign #(in_delay) TIEC440ICURDTOUCHPLBPRIO_delay = TIEC440ICURDTOUCHPLBPRIO;
assign #(in_delay) TIEC440PIR_delay = TIEC440PIR;
assign #(in_delay) TIEC440PVR_delay = TIEC440PVR;
assign #(in_delay) TIEC440USERRESET_delay = TIEC440USERRESET;
assign #(in_delay) TIEDCRBASEADDR_delay = TIEDCRBASEADDR;
assign #(in_delay) TRCC440TRACEDISABLE_delay = TRCC440TRACEDISABLE;
assign #(in_delay) TRCC440TRIGGEREVENTIN_delay = TRCC440TRIGGEREVENTIN;

PPC440_SWIFT ppc440_swift_1 (
	.APU_CONTROL (APU_CONTROL),
	.APU_UDI0 (APU_UDI0),
	.APU_UDI1 (APU_UDI1),
	.APU_UDI10 (APU_UDI10),
	.APU_UDI11 (APU_UDI11),
	.APU_UDI12 (APU_UDI12),
	.APU_UDI13 (APU_UDI13),
	.APU_UDI14 (APU_UDI14),
	.APU_UDI15 (APU_UDI15),
	.APU_UDI2 (APU_UDI2),
	.APU_UDI3 (APU_UDI3),
	.APU_UDI4 (APU_UDI4),
	.APU_UDI5 (APU_UDI5),
	.APU_UDI6 (APU_UDI6),
	.APU_UDI7 (APU_UDI7),
	.APU_UDI8 (APU_UDI8),
	.APU_UDI9 (APU_UDI9),
	.CLOCK_DELAY (CLOCK_DELAY_BINARY),
	.DCR_AUTOLOCK_ENABLE (DCR_AUTOLOCK_ENABLE_BINARY),
	.DMA0_CONTROL (DMA0_CONTROL),
	.DMA0_RXCHANNELCTRL (DMA0_RXCHANNELCTRL),
	.DMA0_RXIRQTIMER (DMA0_RXIRQTIMER),
	.DMA0_TXCHANNELCTRL (DMA0_TXCHANNELCTRL),
	.DMA0_TXIRQTIMER (DMA0_TXIRQTIMER),
	.DMA1_CONTROL (DMA1_CONTROL),
	.DMA1_RXCHANNELCTRL (DMA1_RXCHANNELCTRL),
	.DMA1_RXIRQTIMER (DMA1_RXIRQTIMER),
	.DMA1_TXCHANNELCTRL (DMA1_TXCHANNELCTRL),
	.DMA1_TXIRQTIMER (DMA1_TXIRQTIMER),
	.DMA2_CONTROL (DMA2_CONTROL),
	.DMA2_RXCHANNELCTRL (DMA2_RXCHANNELCTRL),
	.DMA2_RXIRQTIMER (DMA2_RXIRQTIMER),
	.DMA2_TXCHANNELCTRL (DMA2_TXCHANNELCTRL),
	.DMA2_TXIRQTIMER (DMA2_TXIRQTIMER),
	.DMA3_CONTROL (DMA3_CONTROL),
	.DMA3_RXCHANNELCTRL (DMA3_RXCHANNELCTRL),
	.DMA3_RXIRQTIMER (DMA3_RXIRQTIMER),
	.DMA3_TXCHANNELCTRL (DMA3_TXCHANNELCTRL),
	.DMA3_TXIRQTIMER (DMA3_TXIRQTIMER),
	.INTERCONNECT_IMASK (INTERCONNECT_IMASK),
	.INTERCONNECT_TMPL_SEL (INTERCONNECT_TMPL_SEL),
	.MI_ARBCONFIG (MI_ARBCONFIG),
	.MI_BANKCONFLICT_MASK (MI_BANKCONFLICT_MASK),
	.MI_CONTROL (MI_CONTROL),
	.MI_ROWCONFLICT_MASK (MI_ROWCONFLICT_MASK),
	.PPCDM_ASYNCMODE (PPCDM_ASYNCMODE_BINARY),
	.PPCDS_ASYNCMODE (PPCDS_ASYNCMODE_BINARY),
	.PPCM_ARBCONFIG (PPCM_ARBCONFIG),
	.PPCM_CONTROL (PPCM_CONTROL),
	.PPCM_COUNTER (PPCM_COUNTER),
	.PPCS0_ADDRMAP_TMPL0 (PPCS0_ADDRMAP_TMPL0),
	.PPCS0_ADDRMAP_TMPL1 (PPCS0_ADDRMAP_TMPL1),
	.PPCS0_ADDRMAP_TMPL2 (PPCS0_ADDRMAP_TMPL2),
	.PPCS0_ADDRMAP_TMPL3 (PPCS0_ADDRMAP_TMPL3),
	.PPCS0_CONTROL (PPCS0_CONTROL),
	.PPCS0_WIDTH_128N64 (PPCS0_WIDTH_128N64_BINARY),
	.PPCS1_ADDRMAP_TMPL0 (PPCS1_ADDRMAP_TMPL0),
	.PPCS1_ADDRMAP_TMPL1 (PPCS1_ADDRMAP_TMPL1),
	.PPCS1_ADDRMAP_TMPL2 (PPCS1_ADDRMAP_TMPL2),
	.PPCS1_ADDRMAP_TMPL3 (PPCS1_ADDRMAP_TMPL3),
	.PPCS1_CONTROL (PPCS1_CONTROL),
	.PPCS1_WIDTH_128N64 (PPCS1_WIDTH_128N64_BINARY),
	.XBAR_ADDRMAP_TMPL0 (XBAR_ADDRMAP_TMPL0),
	.XBAR_ADDRMAP_TMPL1 (XBAR_ADDRMAP_TMPL1),
	.XBAR_ADDRMAP_TMPL2 (XBAR_ADDRMAP_TMPL2),
	.XBAR_ADDRMAP_TMPL3 (XBAR_ADDRMAP_TMPL3),

	.APUFCMDECFPUOP (APUFCMDECFPUOP_delay),
	.APUFCMDECLDSTXFERSIZE (APUFCMDECLDSTXFERSIZE_delay),
	.APUFCMDECLOAD (APUFCMDECLOAD_delay),
	.APUFCMDECNONAUTON (APUFCMDECNONAUTON_delay),
	.APUFCMDECSTORE (APUFCMDECSTORE_delay),
	.APUFCMDECUDI (APUFCMDECUDI_delay),
	.APUFCMDECUDIVALID (APUFCMDECUDIVALID_delay),
	.APUFCMENDIAN (APUFCMENDIAN_delay),
	.APUFCMFLUSH (APUFCMFLUSH_delay),
	.APUFCMINSTRUCTION (APUFCMINSTRUCTION_delay),
	.APUFCMINSTRVALID (APUFCMINSTRVALID_delay),
	.APUFCMLOADBYTEADDR (APUFCMLOADBYTEADDR_delay),
	.APUFCMLOADDATA (APUFCMLOADDATA_delay),
	.APUFCMLOADDVALID (APUFCMLOADDVALID_delay),
	.APUFCMMSRFE0 (APUFCMMSRFE0_delay),
	.APUFCMMSRFE1 (APUFCMMSRFE1_delay),
	.APUFCMNEXTINSTRREADY (APUFCMNEXTINSTRREADY_delay),
	.APUFCMOPERANDVALID (APUFCMOPERANDVALID_delay),
	.APUFCMRADATA (APUFCMRADATA_delay),
	.APUFCMRBDATA (APUFCMRBDATA_delay),
	.APUFCMWRITEBACKOK (APUFCMWRITEBACKOK_delay),
	.C440CPMCORESLEEPREQ (C440CPMCORESLEEPREQ_delay),
	.C440CPMDECIRPTREQ (C440CPMDECIRPTREQ_delay),
	.C440CPMFITIRPTREQ (C440CPMFITIRPTREQ_delay),
	.C440CPMMSRCE (C440CPMMSRCE_delay),
	.C440CPMMSREE (C440CPMMSREE_delay),
	.C440CPMTIMERRESETREQ (C440CPMTIMERRESETREQ_delay),
	.C440CPMWDIRPTREQ (C440CPMWDIRPTREQ_delay),
	.C440DBGSYSTEMCONTROL (C440DBGSYSTEMCONTROL_delay),
	.C440JTGTDO (C440JTGTDO_delay),
	.C440JTGTDOEN (C440JTGTDOEN_delay),
	.C440MACHINECHECK (C440MACHINECHECK_delay),
	.C440RSTCHIPRESETREQ (C440RSTCHIPRESETREQ_delay),
	.C440RSTCORERESETREQ (C440RSTCORERESETREQ_delay),
	.C440RSTSYSTEMRESETREQ (C440RSTSYSTEMRESETREQ_delay),
	.C440TRCBRANCHSTATUS (C440TRCBRANCHSTATUS_delay),
	.C440TRCCYCLE (C440TRCCYCLE_delay),
	.C440TRCEXECUTIONSTATUS (C440TRCEXECUTIONSTATUS_delay),
	.C440TRCTRACESTATUS (C440TRCTRACESTATUS_delay),
	.C440TRCTRIGGEREVENTOUT (C440TRCTRIGGEREVENTOUT_delay),
	.C440TRCTRIGGEREVENTTYPE (C440TRCTRIGGEREVENTTYPE_delay),
	.DMA0LLRSTENGINEACK (DMA0LLRSTENGINEACK_delay),
	.DMA0LLRXDSTRDYN (DMA0LLRXDSTRDYN_delay),
	.DMA0LLTXD (DMA0LLTXD_delay),
	.DMA0LLTXEOFN (DMA0LLTXEOFN_delay),
	.DMA0LLTXEOPN (DMA0LLTXEOPN_delay),
	.DMA0LLTXREM (DMA0LLTXREM_delay),
	.DMA0LLTXSOFN (DMA0LLTXSOFN_delay),
	.DMA0LLTXSOPN (DMA0LLTXSOPN_delay),
	.DMA0LLTXSRCRDYN (DMA0LLTXSRCRDYN_delay),
	.DMA0RXIRQ (DMA0RXIRQ_delay),
	.DMA0TXIRQ (DMA0TXIRQ_delay),
	.DMA1LLRSTENGINEACK (DMA1LLRSTENGINEACK_delay),
	.DMA1LLRXDSTRDYN (DMA1LLRXDSTRDYN_delay),
	.DMA1LLTXD (DMA1LLTXD_delay),
	.DMA1LLTXEOFN (DMA1LLTXEOFN_delay),
	.DMA1LLTXEOPN (DMA1LLTXEOPN_delay),
	.DMA1LLTXREM (DMA1LLTXREM_delay),
	.DMA1LLTXSOFN (DMA1LLTXSOFN_delay),
	.DMA1LLTXSOPN (DMA1LLTXSOPN_delay),
	.DMA1LLTXSRCRDYN (DMA1LLTXSRCRDYN_delay),
	.DMA1RXIRQ (DMA1RXIRQ_delay),
	.DMA1TXIRQ (DMA1TXIRQ_delay),
	.DMA2LLRSTENGINEACK (DMA2LLRSTENGINEACK_delay),
	.DMA2LLRXDSTRDYN (DMA2LLRXDSTRDYN_delay),
	.DMA2LLTXD (DMA2LLTXD_delay),
	.DMA2LLTXEOFN (DMA2LLTXEOFN_delay),
	.DMA2LLTXEOPN (DMA2LLTXEOPN_delay),
	.DMA2LLTXREM (DMA2LLTXREM_delay),
	.DMA2LLTXSOFN (DMA2LLTXSOFN_delay),
	.DMA2LLTXSOPN (DMA2LLTXSOPN_delay),
	.DMA2LLTXSRCRDYN (DMA2LLTXSRCRDYN_delay),
	.DMA2RXIRQ (DMA2RXIRQ_delay),
	.DMA2TXIRQ (DMA2TXIRQ_delay),
	.DMA3LLRSTENGINEACK (DMA3LLRSTENGINEACK_delay),
	.DMA3LLRXDSTRDYN (DMA3LLRXDSTRDYN_delay),
	.DMA3LLTXD (DMA3LLTXD_delay),
	.DMA3LLTXEOFN (DMA3LLTXEOFN_delay),
	.DMA3LLTXEOPN (DMA3LLTXEOPN_delay),
	.DMA3LLTXREM (DMA3LLTXREM_delay),
	.DMA3LLTXSOFN (DMA3LLTXSOFN_delay),
	.DMA3LLTXSOPN (DMA3LLTXSOPN_delay),
	.DMA3LLTXSRCRDYN (DMA3LLTXSRCRDYN_delay),
	.DMA3RXIRQ (DMA3RXIRQ_delay),
	.DMA3TXIRQ (DMA3TXIRQ_delay),
	.MIMCADDRESS (MIMCADDRESS_delay),
	.MIMCADDRESSVALID (MIMCADDRESSVALID_delay),
	.MIMCBANKCONFLICT (MIMCBANKCONFLICT_delay),
	.MIMCBYTEENABLE (MIMCBYTEENABLE_delay),
	.MIMCREADNOTWRITE (MIMCREADNOTWRITE_delay),
	.MIMCROWCONFLICT (MIMCROWCONFLICT_delay),
	.MIMCWRITEDATA (MIMCWRITEDATA_delay),
	.MIMCWRITEDATAVALID (MIMCWRITEDATAVALID_delay),
	.PPCCPMINTERCONNECTBUSY (PPCCPMINTERCONNECTBUSY_delay),
	.PPCDMDCRABUS (PPCDMDCRABUS_delay),
	.PPCDMDCRDBUSOUT (PPCDMDCRDBUSOUT_delay),
	.PPCDMDCRREAD (PPCDMDCRREAD_delay),
	.PPCDMDCRUABUS (PPCDMDCRUABUS_delay),
	.PPCDMDCRWRITE (PPCDMDCRWRITE_delay),
	.PPCDSDCRACK (PPCDSDCRACK_delay),
	.PPCDSDCRDBUSIN (PPCDSDCRDBUSIN_delay),
	.PPCDSDCRTIMEOUTWAIT (PPCDSDCRTIMEOUTWAIT_delay),
	.PPCEICINTERCONNECTIRQ (PPCEICINTERCONNECTIRQ_delay),
	.PPCMPLBABORT (PPCMPLBABORT_delay),
	.PPCMPLBABUS (PPCMPLBABUS_delay),
	.PPCMPLBBE (PPCMPLBBE_delay),
	.PPCMPLBBUSLOCK (PPCMPLBBUSLOCK_delay),
	.PPCMPLBLOCKERR (PPCMPLBLOCKERR_delay),
	.PPCMPLBPRIORITY (PPCMPLBPRIORITY_delay),
	.PPCMPLBRDBURST (PPCMPLBRDBURST_delay),
	.PPCMPLBREQUEST (PPCMPLBREQUEST_delay),
	.PPCMPLBRNW (PPCMPLBRNW_delay),
	.PPCMPLBSIZE (PPCMPLBSIZE_delay),
	.PPCMPLBTATTRIBUTE (PPCMPLBTATTRIBUTE_delay),
	.PPCMPLBTYPE (PPCMPLBTYPE_delay),
	.PPCMPLBUABUS (PPCMPLBUABUS_delay),
	.PPCMPLBWRBURST (PPCMPLBWRBURST_delay),
	.PPCMPLBWRDBUS (PPCMPLBWRDBUS_delay),
	.PPCS0PLBADDRACK (PPCS0PLBADDRACK_delay),
	.PPCS0PLBMBUSY (PPCS0PLBMBUSY_delay),
	.PPCS0PLBMIRQ (PPCS0PLBMIRQ_delay),
	.PPCS0PLBMRDERR (PPCS0PLBMRDERR_delay),
	.PPCS0PLBMWRERR (PPCS0PLBMWRERR_delay),
	.PPCS0PLBRDBTERM (PPCS0PLBRDBTERM_delay),
	.PPCS0PLBRDCOMP (PPCS0PLBRDCOMP_delay),
	.PPCS0PLBRDDACK (PPCS0PLBRDDACK_delay),
	.PPCS0PLBRDDBUS (PPCS0PLBRDDBUS_delay),
	.PPCS0PLBRDWDADDR (PPCS0PLBRDWDADDR_delay),
	.PPCS0PLBREARBITRATE (PPCS0PLBREARBITRATE_delay),
	.PPCS0PLBSSIZE (PPCS0PLBSSIZE_delay),
	.PPCS0PLBWAIT (PPCS0PLBWAIT_delay),
	.PPCS0PLBWRBTERM (PPCS0PLBWRBTERM_delay),
	.PPCS0PLBWRCOMP (PPCS0PLBWRCOMP_delay),
	.PPCS0PLBWRDACK (PPCS0PLBWRDACK_delay),
	.PPCS1PLBADDRACK (PPCS1PLBADDRACK_delay),
	.PPCS1PLBMBUSY (PPCS1PLBMBUSY_delay),
	.PPCS1PLBMIRQ (PPCS1PLBMIRQ_delay),
	.PPCS1PLBMRDERR (PPCS1PLBMRDERR_delay),
	.PPCS1PLBMWRERR (PPCS1PLBMWRERR_delay),
	.PPCS1PLBRDBTERM (PPCS1PLBRDBTERM_delay),
	.PPCS1PLBRDCOMP (PPCS1PLBRDCOMP_delay),
	.PPCS1PLBRDDACK (PPCS1PLBRDDACK_delay),
	.PPCS1PLBRDDBUS (PPCS1PLBRDDBUS_delay),
	.PPCS1PLBRDWDADDR (PPCS1PLBRDWDADDR_delay),
	.PPCS1PLBREARBITRATE (PPCS1PLBREARBITRATE_delay),
	.PPCS1PLBSSIZE (PPCS1PLBSSIZE_delay),
	.PPCS1PLBWAIT (PPCS1PLBWAIT_delay),
	.PPCS1PLBWRBTERM (PPCS1PLBWRBTERM_delay),
	.PPCS1PLBWRCOMP (PPCS1PLBWRCOMP_delay),
	.PPCS1PLBWRDACK (PPCS1PLBWRDACK_delay),

	.CPMC440CLK (CPMC440CLK_delay),
	.CPMC440CLKEN (CPMC440CLKEN_delay),
	.CPMC440CORECLOCKINACTIVE (CPMC440CORECLOCKINACTIVE_delay),
	.CPMC440TIMERCLOCK (CPMC440TIMERCLOCK_delay),
	.CPMDCRCLK (CPMDCRCLK_delay),
	.CPMDMA0LLCLK (CPMDMA0LLCLK_delay),
	.CPMDMA1LLCLK (CPMDMA1LLCLK_delay),
	.CPMDMA2LLCLK (CPMDMA2LLCLK_delay),
	.CPMDMA3LLCLK (CPMDMA3LLCLK_delay),
	.CPMFCMCLK (CPMFCMCLK_delay),
	.CPMINTERCONNECTCLK (CPMINTERCONNECTCLK_delay),
	.CPMINTERCONNECTCLKEN (CPMINTERCONNECTCLKEN_delay),
	.CPMINTERCONNECTCLKNTO1 (CPMINTERCONNECTCLKNTO1_delay),
	.CPMMCCLK (CPMMCCLK_delay),
	.CPMPPCMPLBCLK (CPMPPCMPLBCLK_delay),
	.CPMPPCS0PLBCLK (CPMPPCS0PLBCLK_delay),
	.CPMPPCS1PLBCLK (CPMPPCS1PLBCLK_delay),
	.DBGC440DEBUGHALT (DBGC440DEBUGHALT_delay),
	.DBGC440SYSTEMSTATUS (DBGC440SYSTEMSTATUS_delay),
	.DBGC440UNCONDDEBUGEVENT (DBGC440UNCONDDEBUGEVENT_delay),
	.DCRPPCDMACK (DCRPPCDMACK_delay),
	.DCRPPCDMDBUSIN (DCRPPCDMDBUSIN_delay),
	.DCRPPCDMTIMEOUTWAIT (DCRPPCDMTIMEOUTWAIT_delay),
	.DCRPPCDSABUS (DCRPPCDSABUS_delay),
	.DCRPPCDSDBUSOUT (DCRPPCDSDBUSOUT_delay),
	.DCRPPCDSREAD (DCRPPCDSREAD_delay),
	.DCRPPCDSWRITE (DCRPPCDSWRITE_delay),
	.EICC440CRITIRQ (EICC440CRITIRQ_delay),
	.EICC440EXTIRQ (EICC440EXTIRQ_delay),
	.FCMAPUCONFIRMINSTR (FCMAPUCONFIRMINSTR_delay),
	.FCMAPUCR (FCMAPUCR_delay),
	.FCMAPUDONE (FCMAPUDONE_delay),
	.FCMAPUEXCEPTION (FCMAPUEXCEPTION_delay),
	.FCMAPUFPSCRFEX (FCMAPUFPSCRFEX_delay),
	.FCMAPURESULT (FCMAPURESULT_delay),
	.FCMAPURESULTVALID (FCMAPURESULTVALID_delay),
	.FCMAPUSLEEPNOTREADY (FCMAPUSLEEPNOTREADY_delay),
	.FCMAPUSTOREDATA (FCMAPUSTOREDATA_delay),
	.JTGC440TCK (JTGC440TCK_delay),
	.JTGC440TDI (JTGC440TDI_delay),
	.JTGC440TMS (JTGC440TMS_delay),
	.JTGC440TRSTNEG (JTGC440TRSTNEG_delay),
	.LLDMA0RSTENGINEREQ (LLDMA0RSTENGINEREQ_delay),
	.LLDMA0RXD (LLDMA0RXD_delay),
	.LLDMA0RXEOFN (LLDMA0RXEOFN_delay),
	.LLDMA0RXEOPN (LLDMA0RXEOPN_delay),
	.LLDMA0RXREM (LLDMA0RXREM_delay),
	.LLDMA0RXSOFN (LLDMA0RXSOFN_delay),
	.LLDMA0RXSOPN (LLDMA0RXSOPN_delay),
	.LLDMA0RXSRCRDYN (LLDMA0RXSRCRDYN_delay),
	.LLDMA0TXDSTRDYN (LLDMA0TXDSTRDYN_delay),
	.LLDMA1RSTENGINEREQ (LLDMA1RSTENGINEREQ_delay),
	.LLDMA1RXD (LLDMA1RXD_delay),
	.LLDMA1RXEOFN (LLDMA1RXEOFN_delay),
	.LLDMA1RXEOPN (LLDMA1RXEOPN_delay),
	.LLDMA1RXREM (LLDMA1RXREM_delay),
	.LLDMA1RXSOFN (LLDMA1RXSOFN_delay),
	.LLDMA1RXSOPN (LLDMA1RXSOPN_delay),
	.LLDMA1RXSRCRDYN (LLDMA1RXSRCRDYN_delay),
	.LLDMA1TXDSTRDYN (LLDMA1TXDSTRDYN_delay),
	.LLDMA2RSTENGINEREQ (LLDMA2RSTENGINEREQ_delay),
	.LLDMA2RXD (LLDMA2RXD_delay),
	.LLDMA2RXEOFN (LLDMA2RXEOFN_delay),
	.LLDMA2RXEOPN (LLDMA2RXEOPN_delay),
	.LLDMA2RXREM (LLDMA2RXREM_delay),
	.LLDMA2RXSOFN (LLDMA2RXSOFN_delay),
	.LLDMA2RXSOPN (LLDMA2RXSOPN_delay),
	.LLDMA2RXSRCRDYN (LLDMA2RXSRCRDYN_delay),
	.LLDMA2TXDSTRDYN (LLDMA2TXDSTRDYN_delay),
	.LLDMA3RSTENGINEREQ (LLDMA3RSTENGINEREQ_delay),
	.LLDMA3RXD (LLDMA3RXD_delay),
	.LLDMA3RXEOFN (LLDMA3RXEOFN_delay),
	.LLDMA3RXEOPN (LLDMA3RXEOPN_delay),
	.LLDMA3RXREM (LLDMA3RXREM_delay),
	.LLDMA3RXSOFN (LLDMA3RXSOFN_delay),
	.LLDMA3RXSOPN (LLDMA3RXSOPN_delay),
	.LLDMA3RXSRCRDYN (LLDMA3RXSRCRDYN_delay),
	.LLDMA3TXDSTRDYN (LLDMA3TXDSTRDYN_delay),
	.MCMIADDRREADYTOACCEPT (MCMIADDRREADYTOACCEPT_delay),
	.MCMIREADDATA (MCMIREADDATA_delay),
	.MCMIREADDATAERR (MCMIREADDATAERR_delay),
	.MCMIREADDATAVALID (MCMIREADDATAVALID_delay),
	.PLBPPCMADDRACK (PLBPPCMADDRACK_delay),
	.PLBPPCMMBUSY (PLBPPCMMBUSY_delay),
	.PLBPPCMMIRQ (PLBPPCMMIRQ_delay),
	.PLBPPCMMRDERR (PLBPPCMMRDERR_delay),
	.PLBPPCMMWRERR (PLBPPCMMWRERR_delay),
	.PLBPPCMRDBTERM (PLBPPCMRDBTERM_delay),
	.PLBPPCMRDDACK (PLBPPCMRDDACK_delay),
	.PLBPPCMRDDBUS (PLBPPCMRDDBUS_delay),
	.PLBPPCMRDPENDPRI (PLBPPCMRDPENDPRI_delay),
	.PLBPPCMRDPENDREQ (PLBPPCMRDPENDREQ_delay),
	.PLBPPCMRDWDADDR (PLBPPCMRDWDADDR_delay),
	.PLBPPCMREARBITRATE (PLBPPCMREARBITRATE_delay),
	.PLBPPCMREQPRI (PLBPPCMREQPRI_delay),
	.PLBPPCMSSIZE (PLBPPCMSSIZE_delay),
	.PLBPPCMTIMEOUT (PLBPPCMTIMEOUT_delay),
	.PLBPPCMWRBTERM (PLBPPCMWRBTERM_delay),
	.PLBPPCMWRDACK (PLBPPCMWRDACK_delay),
	.PLBPPCMWRPENDPRI (PLBPPCMWRPENDPRI_delay),
	.PLBPPCMWRPENDREQ (PLBPPCMWRPENDREQ_delay),
	.PLBPPCS0ABORT (PLBPPCS0ABORT_delay),
	.PLBPPCS0ABUS (PLBPPCS0ABUS_delay),
	.PLBPPCS0BE (PLBPPCS0BE_delay),
	.PLBPPCS0BUSLOCK (PLBPPCS0BUSLOCK_delay),
	.PLBPPCS0LOCKERR (PLBPPCS0LOCKERR_delay),
	.PLBPPCS0MASTERID (PLBPPCS0MASTERID_delay),
	.PLBPPCS0MSIZE (PLBPPCS0MSIZE_delay),
	.PLBPPCS0PAVALID (PLBPPCS0PAVALID_delay),
	.PLBPPCS0RDBURST (PLBPPCS0RDBURST_delay),
	.PLBPPCS0RDPENDPRI (PLBPPCS0RDPENDPRI_delay),
	.PLBPPCS0RDPENDREQ (PLBPPCS0RDPENDREQ_delay),
	.PLBPPCS0RDPRIM (PLBPPCS0RDPRIM_delay),
	.PLBPPCS0REQPRI (PLBPPCS0REQPRI_delay),
	.PLBPPCS0RNW (PLBPPCS0RNW_delay),
	.PLBPPCS0SAVALID (PLBPPCS0SAVALID_delay),
	.PLBPPCS0SIZE (PLBPPCS0SIZE_delay),
	.PLBPPCS0TATTRIBUTE (PLBPPCS0TATTRIBUTE_delay),
	.PLBPPCS0TYPE (PLBPPCS0TYPE_delay),
	.PLBPPCS0UABUS (PLBPPCS0UABUS_delay),
	.PLBPPCS0WRBURST (PLBPPCS0WRBURST_delay),
	.PLBPPCS0WRDBUS (PLBPPCS0WRDBUS_delay),
	.PLBPPCS0WRPENDPRI (PLBPPCS0WRPENDPRI_delay),
	.PLBPPCS0WRPENDREQ (PLBPPCS0WRPENDREQ_delay),
	.PLBPPCS0WRPRIM (PLBPPCS0WRPRIM_delay),
	.PLBPPCS1ABORT (PLBPPCS1ABORT_delay),
	.PLBPPCS1ABUS (PLBPPCS1ABUS_delay),
	.PLBPPCS1BE (PLBPPCS1BE_delay),
	.PLBPPCS1BUSLOCK (PLBPPCS1BUSLOCK_delay),
	.PLBPPCS1LOCKERR (PLBPPCS1LOCKERR_delay),
	.PLBPPCS1MASTERID (PLBPPCS1MASTERID_delay),
	.PLBPPCS1MSIZE (PLBPPCS1MSIZE_delay),
	.PLBPPCS1PAVALID (PLBPPCS1PAVALID_delay),
	.PLBPPCS1RDBURST (PLBPPCS1RDBURST_delay),
	.PLBPPCS1RDPENDPRI (PLBPPCS1RDPENDPRI_delay),
	.PLBPPCS1RDPENDREQ (PLBPPCS1RDPENDREQ_delay),
	.PLBPPCS1RDPRIM (PLBPPCS1RDPRIM_delay),
	.PLBPPCS1REQPRI (PLBPPCS1REQPRI_delay),
	.PLBPPCS1RNW (PLBPPCS1RNW_delay),
	.PLBPPCS1SAVALID (PLBPPCS1SAVALID_delay),
	.PLBPPCS1SIZE (PLBPPCS1SIZE_delay),
	.PLBPPCS1TATTRIBUTE (PLBPPCS1TATTRIBUTE_delay),
	.PLBPPCS1TYPE (PLBPPCS1TYPE_delay),
	.PLBPPCS1UABUS (PLBPPCS1UABUS_delay),
	.PLBPPCS1WRBURST (PLBPPCS1WRBURST_delay),
	.PLBPPCS1WRDBUS (PLBPPCS1WRDBUS_delay),
	.PLBPPCS1WRPENDPRI (PLBPPCS1WRPENDPRI_delay),
	.PLBPPCS1WRPENDREQ (PLBPPCS1WRPENDREQ_delay),
	.PLBPPCS1WRPRIM (PLBPPCS1WRPRIM_delay),
	.RSTC440RESETCHIP (RSTC440RESETCHIP_delay),
	.RSTC440RESETCORE (RSTC440RESETCORE_delay),
	.RSTC440RESETSYSTEM (RSTC440RESETSYSTEM_delay),
	.TIEC440DCURDLDCACHEPLBPRIO (TIEC440DCURDLDCACHEPLBPRIO_delay),
	.TIEC440DCURDNONCACHEPLBPRIO (TIEC440DCURDNONCACHEPLBPRIO_delay),
	.TIEC440DCURDTOUCHPLBPRIO (TIEC440DCURDTOUCHPLBPRIO_delay),
	.TIEC440DCURDURGENTPLBPRIO (TIEC440DCURDURGENTPLBPRIO_delay),
	.TIEC440DCUWRFLUSHPLBPRIO (TIEC440DCUWRFLUSHPLBPRIO_delay),
	.TIEC440DCUWRSTOREPLBPRIO (TIEC440DCUWRSTOREPLBPRIO_delay),
	.TIEC440DCUWRURGENTPLBPRIO (TIEC440DCUWRURGENTPLBPRIO_delay),
	.TIEC440ENDIANRESET (TIEC440ENDIANRESET_delay),
	.TIEC440ERPNRESET (TIEC440ERPNRESET_delay),
	.TIEC440ICURDFETCHPLBPRIO (TIEC440ICURDFETCHPLBPRIO_delay),
	.TIEC440ICURDSPECPLBPRIO (TIEC440ICURDSPECPLBPRIO_delay),
	.TIEC440ICURDTOUCHPLBPRIO (TIEC440ICURDTOUCHPLBPRIO_delay),
	.TIEC440PIR (TIEC440PIR_delay),
	.TIEC440PVR (TIEC440PVR_delay),
	.TIEC440USERRESET (TIEC440USERRESET_delay),
	.TIEDCRBASEADDR (TIEDCRBASEADDR_delay),
	.TRCC440TRACEDISABLE (TRCC440TRACEDISABLE_delay),
	.TRCC440TRIGGEREVENTIN (TRCC440TRIGGEREVENTIN_delay),
	.GSR (GSR)
);

specify
	(CPMC440CLK => C440CPMCORESLEEPREQ) = (100, 100);
	(CPMC440CLK => C440CPMDECIRPTREQ) = (100, 100);
	(CPMC440CLK => C440CPMFITIRPTREQ) = (100, 100);
	(CPMC440CLK => C440CPMMSRCE) = (100, 100);
	(CPMC440CLK => C440CPMMSREE) = (100, 100);
	(CPMC440CLK => C440CPMTIMERRESETREQ) = (100, 100);
	(CPMC440CLK => C440CPMWDIRPTREQ) = (100, 100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL) = (100, 100);
	(CPMC440CLK => C440MACHINECHECK) = (100, 100);
	(CPMC440CLK => C440TRCBRANCHSTATUS) = (100, 100);
	(CPMC440CLK => C440TRCCYCLE) = (100, 100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS) = (100, 100);
	(CPMC440CLK => C440TRCTRACESTATUS) = (100, 100);
	(CPMC440CLK => C440TRCTRIGGEREVENTOUT) = (100, 100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE) = (100, 100);
	(CPMDCRCLK => PPCDMDCRABUS) = (100, 100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT) = (100, 100);
	(CPMDCRCLK => PPCDMDCRREAD) = (100, 100);
	(CPMDCRCLK => PPCDMDCRUABUS) = (100, 100);
	(CPMDCRCLK => PPCDMDCRWRITE) = (100, 100);
	(CPMDCRCLK => PPCDSDCRACK) = (100, 100);
	(CPMDCRCLK => PPCDSDCRDBUSIN) = (100, 100);
	(CPMDCRCLK => PPCDSDCRTIMEOUTWAIT) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLRSTENGINEACK) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLRXDSTRDYN) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXD) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXEOFN) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXEOPN) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXREM) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXSOFN) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXSOPN) = (100, 100);
	(CPMDMA0LLCLK => DMA0LLTXSRCRDYN) = (100, 100);
	(CPMDMA0LLCLK => DMA0RXIRQ) = (100, 100);
	(CPMDMA0LLCLK => DMA0TXIRQ) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLRSTENGINEACK) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLRXDSTRDYN) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXD) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXEOFN) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXEOPN) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXREM) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXSOFN) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXSOPN) = (100, 100);
	(CPMDMA1LLCLK => DMA1LLTXSRCRDYN) = (100, 100);
	(CPMDMA1LLCLK => DMA1RXIRQ) = (100, 100);
	(CPMDMA1LLCLK => DMA1TXIRQ) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLRSTENGINEACK) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLRXDSTRDYN) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXD) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXEOFN) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXEOPN) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXREM) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXSOFN) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXSOPN) = (100, 100);
	(CPMDMA2LLCLK => DMA2LLTXSRCRDYN) = (100, 100);
	(CPMDMA2LLCLK => DMA2RXIRQ) = (100, 100);
	(CPMDMA2LLCLK => DMA2TXIRQ) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLRSTENGINEACK) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLRXDSTRDYN) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXD) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXEOFN) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXEOPN) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXREM) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXSOFN) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXSOPN) = (100, 100);
	(CPMDMA3LLCLK => DMA3LLTXSRCRDYN) = (100, 100);
	(CPMDMA3LLCLK => DMA3RXIRQ) = (100, 100);
	(CPMDMA3LLCLK => DMA3TXIRQ) = (100, 100);
	(CPMFCMCLK => APUFCMDECFPUOP) = (100, 100);
	(CPMFCMCLK => APUFCMDECLDSTXFERSIZE) = (100, 100);
	(CPMFCMCLK => APUFCMDECLOAD) = (100, 100);
	(CPMFCMCLK => APUFCMDECNONAUTON) = (100, 100);
	(CPMFCMCLK => APUFCMDECSTORE) = (100, 100);
	(CPMFCMCLK => APUFCMDECUDI) = (100, 100);
	(CPMFCMCLK => APUFCMDECUDIVALID) = (100, 100);
	(CPMFCMCLK => APUFCMENDIAN) = (100, 100);
	(CPMFCMCLK => APUFCMFLUSH) = (100, 100);
	(CPMFCMCLK => APUFCMINSTRUCTION) = (100, 100);
	(CPMFCMCLK => APUFCMINSTRVALID) = (100, 100);
	(CPMFCMCLK => APUFCMLOADBYTEADDR) = (100, 100);
	(CPMFCMCLK => APUFCMLOADDATA) = (100, 100);
	(CPMFCMCLK => APUFCMLOADDVALID) = (100, 100);
	(CPMFCMCLK => APUFCMMSRFE0) = (100, 100);
	(CPMFCMCLK => APUFCMMSRFE1) = (100, 100);
	(CPMFCMCLK => APUFCMNEXTINSTRREADY) = (100, 100);
	(CPMFCMCLK => APUFCMOPERANDVALID) = (100, 100);
	(CPMFCMCLK => APUFCMRADATA) = (100, 100);
	(CPMFCMCLK => APUFCMRBDATA) = (100, 100);
	(CPMFCMCLK => APUFCMWRITEBACKOK) = (100, 100);
	(CPMINTERCONNECTCLK => C440RSTCHIPRESETREQ) = (100, 100);
	(CPMINTERCONNECTCLK => C440RSTCORERESETREQ) = (100, 100);
	(CPMINTERCONNECTCLK => C440RSTSYSTEMRESETREQ) = (100, 100);
	(CPMINTERCONNECTCLK => PPCCPMINTERCONNECTBUSY) = (100, 100);
	(CPMINTERCONNECTCLK => PPCEICINTERCONNECTIRQ) = (100, 100);
	(CPMMCCLK => MIMCADDRESS) = (100, 100);
	(CPMMCCLK => MIMCADDRESSVALID) = (100, 100);
	(CPMMCCLK => MIMCBANKCONFLICT) = (100, 100);
	(CPMMCCLK => MIMCBYTEENABLE) = (100, 100);
	(CPMMCCLK => MIMCREADNOTWRITE) = (100, 100);
	(CPMMCCLK => MIMCROWCONFLICT) = (100, 100);
	(CPMMCCLK => MIMCWRITEDATA) = (100, 100);
	(CPMMCCLK => MIMCWRITEDATAVALID) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBABORT) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBABUS) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBBE) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBBUSLOCK) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBLOCKERR) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBPRIORITY) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBRDBURST) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBREQUEST) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBRNW) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBSIZE) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBTYPE) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBUABUS) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBWRBURST) = (100, 100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBADDRACK) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBMBUSY) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBMIRQ) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBMRDERR) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBMWRERR) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDBTERM) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDCOMP) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDACK) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDWDADDR) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBREARBITRATE) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBSSIZE) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBWAIT) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRBTERM) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRCOMP) = (100, 100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRDACK) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBADDRACK) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBMBUSY) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBMIRQ) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBMRDERR) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBMWRERR) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDBTERM) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDCOMP) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDACK) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDWDADDR) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBREARBITRATE) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBSSIZE) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBWAIT) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRBTERM) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRCOMP) = (100, 100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRDACK) = (100, 100);
	(JTGC440TCK => C440JTGTDO) = (100, 100);
	(JTGC440TCK => C440JTGTDOEN) = (100, 100);
	specparam PATHPULSE$ = 0;
endspecify
endmodule
